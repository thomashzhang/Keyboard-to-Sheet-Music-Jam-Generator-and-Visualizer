BZh91AY&SY�N�,��߀pp���f� ?���a|� (z!
!A%�TE*�RB�J$�P��
�I!%R��R�I��>��$P �@      %
(������ �Q$� "���J��P��*H���   ��   $
 �8�t �$��������` �t��=��tr�{n��졛|A�� N!��&���w��s��;��\�v�S��ZV�t��{� �T�b{j�n���m�V��9��@
Q�j��  P    V�tv;ݫ*qn��Ys3����@=�K>��iye��W���J^� �K;=�G�W  = �l.m�5]� {�Qr{��FJ�Uv�^�_zT�T�[����\�_crj��� � 
   c� ��Q��.6\c\ڥ��׳�� �s��&�Nm�C�y�*��ek� ��������t�  W�UK=��ϥ <�cIYe�Vs�N�MɻZۀF�{5�7���g����c�ݛg&� {��   ( ��>>�>��7L�i]��U{���
7�I\�|��x�{4��g�x�KA@里��2��8  ���Y��^<} �<�+-�gG�ݍťS{��@���ڎ{8����g�:�� ��P ( %��P���st�F|cqa�9�z<��*'y���>�w��o�Ey���<�  c��ۛR=� �Tc>��C�W�g�wk�������OW��<��3��8P       ��ةJ��` �y&& 4��CR����zL���'�UJ�  Ѡ    D�*���$�`�4�0&	������MT�UF� �4b R%(��Dȣ�OS#@h�jfS�O���_�/������{{}�^�QTUW���B����PUT�R������Ȩ���#i�M���?���EUkUEU{��/�!UW��t������U���������/�X���[kV/�gS��^�+Y��?�Ȩ�5��kX%.�4u�3Y��	BP�2g{
��^��8��W+)�-Vʾ6�:+�y�y@�E �:�JN��;=؅Eh�
6�
$��ŧx&Q�][taq!9�/x�\Dm5�װ{u�%I��]V,a�r	:����>U��Д7N�	�K����vu'�Ã�Nןi�����-�Z��w	���u�zd�k]��<��F�J�L�j�]���꥕���<�n-H�s��pQv�B6Sn�@S��Mg�Buj�˜����s�"�MS:#��)	�K(��e�̟ǻGn�E��V�vm۽��>�w�5<B�GV�r/y���\ T��9�XY��绢�q{%^P���V5b�9|Ǔ�v+M�S�X*@�}��Ʊ�?zq�R����)4u�x�wbll��aJR�iX Bj�I��y�S�xM^Z~��܀��F��J�Q��5�SA�PK��s0��Iubh����*)z�r�X`�麵��a��D +i�Qe�)Z�{՜8�K�b�Z*A]��Z98V-j�R��L���*��0��l�%�Æ���upm�iΩb�bey,��\G��Q�.�!,E�(��DK[�����f���mj*n�&�5���rLxj���Ѳ��F��h���rx����AD�Z5�����tbZ81&բ��w���Iv���G��%	�;7���h�a�볨N��'Z��u�����ģu�DHg7�Ө�j͛�f=�=���^�ו�º��;Ӕ�LMB�`�G�йC�2��*��ubH1jBLThZ��V���uq��|�F�/����;����Xq�0��:MK��	�C�Q�;�Ðb�&�-9޿^
qC�U�E	�j���W���d�8�����Y5TZՂ��ڈb���N��ļ�'�N��UΕ��TW�Zؐ�fu�x�����w�]8^RbK�����(;����;(�w	��&�oo5���'�j#!�fd�%ȣ�ȍy޺�5����6���t����ļY�ֻǈR���!X��z�'YTcFQ׃�y����C��N�|�\�հ&մ�:B����Y�)ɔ <�u��t�Z�z��^��|�L�*ok� ���j݉K�&DY���Mk{���2�2)ők@��_x�\9Qu崢�AR�]b��~���O�.��	��6�e�z�#Q��X�tZ�S$�v�"01���qc�=�.-��d��tw�х�eǣa�	[s��`�ԚL�GON���k0'��0����:]X���]�W��گV��BP�%	�'����{�F��{�\�M�ƉHb9w:.
��`{h+7�ׁ���	BP��nP�	�N�8Bn��(J�J��M�&�7	�N�5	�%	Bu�P���z%�q����k/tg�{��^�y�����,\jע��K�W\]B�P���*�����%�YU�5yl��k���ͷցp�K:�w\B���ӥmx�=a��Q�2u���U)/$�tJηW\���F.)q�H�a'Ŋ��Р�s]WD�w��]V��+�*��ȵ:�����F��(�l�ך�ӨOa2]��5��Br�q�Ju���15j���M��li��2��t<�V��j�|���9�궔�MZ�p]%�ЉY��ƫ�t�������������*�*��К;��F5��%� �F�JPY���mkk�5�VN׌��k;�J39iN����/No/6
�r��V����X��a��u��:�)��z6�9kHd�$�b��Ɗ�W�Ӫvع�'q �&�z����]m���(J��-ë3��c���6p<�k��Z�j�����)o2�{��xW��JȲ׺��n�[m.īcT�*F+X�ۡ9��<�]��G�6�# ��{�a�J��9�{4�n�j�Q��lnm�l�Z��*@���(MBP�%�S���ىw�S����C���l�jٞ�1,+����Q<�vr��,/
��T���(J_u���i��D��3go�&BP�	BP�RH){�H���P��ֵ~Ą[X��Q�f
q�W�xK����Ư�����7��|�Rԗ��5UR�=��R��!�(���^K����,�.��&�D�A<hۄf]p;�y�:�{�.�v�r�[)[�J��O���U��J'VD,�<N�����~juN�b�⒞��:���8��&�w�s]���ý�s�h-5����Ü����]Qw��r�+]�_&#'pF�@���L��#��<���a�E,�j4A�r�X)���N�vZ�H¼��;��:�)�%-�BVŔݠMq.\}Ga䳉X�\F��Bo1	�:��(�Ks��)]	yb�
�&�l'j�'e3���yA+�|Ev]��IdK�mp��K��*e$�L�_gu%b�p�'��H{���;#<����vo��p���29���y�20��Ӻd罛o��yR�HLe
�K��v�
���/�.	:玘�I�.WW$�Y��k�ӡ������ �K1���P�%���!6�̎�w�p�p�~��P�;dO������Q"��R���\MNv�|K!pRTMuu:�J�YY��V�Ǧ��E&Q�3}GK�K���.��s&�V0o��t�Åc��ᳳ�lÎ��Od�P]��"L�c�Ԛ����o���BP������;��&�(MBj|z��F�y�w��pyc�F�uؔ&�2�{���ѷ:jWD��dR���Z�-L�/5!�v���łiy<�ӓ�Γ�ޝB睤&��.��̮'�<��\w)Ҽ�|�2����^�.VuI�ib�*@�u�KH]��y�z�Z����F��5�n��&˯y�t9a�qq���'(W|��=��1�3�t���ٜ�l�V*Xڥ�RHu��l[j��.N�1��v����乍Z����4�\*(�j�LB[��qF�U��l#����8��DՕ'x㤤�)�v�
!(NBP��P�=���;;234l2�r����\�P��`�/5&6�Mk��j�ā "�DTNdw�G��J!=��������i�E;4�]94T�7'I�����\<�BP�%�֌�+��h�M�̈��	�yk�p��me8uQky�Uu�鼃[5�l��=!(JR�0r��ч[�5��ٱ���r�Y"IC��ܝ�e�z��如���,A�eLT���v�%G �Nv&f��Q��)�߶�
����E����9���qu������r��Ҕ��H�YJ�cI�-�Y��<�P�%)�y��4h���[�U�'V�\�V&���v�R�R
�ZGJ(�*���7��<��L���B�+��k�̊�ӫ�9��Ug ����b}]uuW�[c�Zʺ����f�]���C�Y�/^�S��m:�W>�F]Zb�;�!;��'$7�{���PĘ����<)]�RitN����������Mb�G(�M+�N�QbĊ��C��N�PR WlR YK��Z�z	5j.��*q�:��7��dx�;w-�Y�q;�.������Æ����
&4�99���H�Y�E���5��{�3j�4��DE��y��4J�唑�8���Sk՗�u�N��	���+r�<����]<Sq>���q.dt�m;h��0��EJ
�(�bAC�+Qo.�x��*���1u����%	���u	BjSp�p���zt�k��v��3�bV��x%"\B���%�yz��N{��"�SuӽN�3�款�@�P���X���:���P�Yd�YI�`F`��4�0�V5䅑	�������v��eqV�H/`v�$��Q���pE�ibE��S�*�H.WJvJ�o=�]z�e�k9�{'11ǧq#�gS�Rw-C9�vgl�!֋Q�d�N���`ԙ�h��f!�:`�34G}�J�ί\R���W:�YN�İ\Υ���&�@Pt����ıB���S7��'V�C�:}cV��v�����$ڲ�PE�ڡX���VV
�g�+WӨ1ۨċ%ӒF�ֳ\�ܵtNQ�
9LI�b � oN���D+Qp�$�%�EI����m�9�'����3 ��ʡ;�ή�R��YK�V`��v��&<K��/X��<�Z��-\̑=��|�V��Qw��][W�r�JOy4��"3 ԙ�4�77Y�3Wv�Qʳ8:�.�B���y�������v�yA��Yt�(�y(�(��T�܎�^*�w�bf>���K6p�]�����9at:�N�&����[�]�W���w��u�<.U]�Q�F�u�r4V���{	���9(�;�Yj�S�����qE�%�����p�u�W8'9#S���:�j<��( 7���;��y�����T�Z��k��;}���V��:����V5u���w�k��m]���\���N����^O��8RUY��&�]Ψ�ܮ���j�/����b�uq�
+*I��9�f�Wt��;��N{���s�Rd�牉�c�5h�xi��εю�Ԙ�	biYV2�V��Y\\Q���&($�0���]8��\K
��(�U��ST93Ej\sC�dc��8I��A�y���w#�Zua0e�ju���a:J΢��W�Dr�_;����]q��S V�j�#��C\3؍��cP�A�]��R�X(�E+�.VQm:��Pdh���7dkB��kM��������%�����"P��HCv�/��o���\C!)�	�����vSκPK��P�R�y2����X��b��Н��Q�ѿF��%� ��Z7.��\��U���'`�Յ���I%TUe�������uo�:p|׌a������ym��	�k#Qfj�fuGy���]=A�j|�ӑ�{�a�{[�O�����i�kxN:�0�q�[xow�P�&Hk4�9�{��GI�K�j۠-	t/)�喕�p~t(��S�.��R�:�R'-�W{i[��,E>w�����Խ��9X���Ӥ�wmzw[
�/-Wl��f�c�Em�tX�Y���
��u2�R;�e�#ɶ����   8    v�            C�    �                   m�           9oZ�sM���ml��l nu�&Iev�]���pM�`�E���g����j۶�Vr=�C³�k�� 6���j��z�m�Ѯ�M�I  �llYv�j�L���|��cgk�P��M�1�X��=��������xT��Ağ7�i>כm������k f��6�`Ut!6�Rpn�R6ݺ8�1��<��P�s�m�~|6�*�_�ƻm����CQ�q����*R۶.$	X�m�L;f�ZD{M�Ҡ5���#�i��-��u0�Mb2'Z���z]��*��][d�3��ɒ��R٘祐*�Ir���MX�%T�X��{L�UW:إ�&e69�B��		���u���:CM����J���t��U<�J�t�Κ� �Cm���l�%��$6k�ݫ�ؠ�q���(幄d�j�]��N��    ���` p�|    z�      h   �l      $                                    ��(0 8��  �J �@
Pan�  6�      >>��    �8            Y@             ��    ׭              %�     �>  8 �      �(    �    �i6	     3�   �  ���        � C sE"�
Q���  �$p (0� �P`8 p +� �   �����l�   8 p +�lA�����!���0 8����)@A��߶���w�  $� �p	     � $    ��   K���.�`�o�ŷ��klQ���k�B�=��]UW5)'NZ/�n[wmr�u�L�t�F    I���Ͷݱ'�],ԫ]R*�c@枝]��< &��kg��l���[���4+f���C"���]"�.�H�7q�� Ù[WY���^y�j��;�v���A��e��jK�z*�Y;k�.��ʽ�ɨ�MJ:��-�6�m�kX-幀��DȺ��Z�U
�UU^�{GB��[��`]*�FCv��cz�v��ւ�2$�R��zN���X�f����T�7��{`��	B���T�ę-rg�E��qWl�@Q�UUA�<'A�6I�͎K��ǪW��v����r))�;v�+���SԎ�^�'.�AV:rK���(1)yg�j��z�Wg��V��5�X�ٶr���re��Uml���.,�M�ѹPiԭ�U:ز��-�$����
�mCS����x^�bu�-�왙��6�L!�U۳-��㬄�[L�Qq3tjy]�p�u�(J���[�/��a X�n�!su�X6ت��鬀��v�q�ԣ�"m���ܾd�"36��L2�o$t�{3R���j���g�l��P ��$*sp��E�9��:�u�g/JI&�;l���Ď7i���h �^�I�����)v[r��}o����]$PJ�vTȪ�+5UmR�Us���RW��Iw�-�h<d^�`���6�@ID�UU��ث[�ۅ��)�ɑU�t��1��z@�D��R�d��|���i�6��-%���q���f�T��3*���HYF�+<͊ Xy�����]�-�:vt��֒���X�Qg5PB�X-��UV�PZ��y�*�E]�m��P���@:\�{f�@ �6݇^۱�)���BMLʄ:{g�`�Bj�#R�]i9�KnQ֌�7l���� �*e�Ĳ��V�ۂ.:i�]��V�fD�m�pٳl-6�7V�[@ ��!s[���X��ə�avW�����b&���[iVVykְmUյclU��	�kj���E�iybܓ�T=�K���6�� [7E�(�6����+(UT�qJ��9,��#[*���/FR����Ɛ6�� �n��l����h2Kd��t��А��ր:��k"�V��эZ���P�x�S�8"UkSh�j��iV�꫁�����d���FIj����U�j��
�hhδnA@�z$;,��ngk��9Q�8�q�˴�h*���*�WW7-!;x�L��R��k��������ı��K+��WT�\���\k�z���+J���v��YWHV�um*�U�;t��(|�� �Eχ;?.�Q��d.hD���@�VN�ʱ�����
L��HZ3j�ä�x��[@5�@횧B�*�UUT�*�Y%.@v�Z��qh�-��6�m��T��8�U�Mn��l�ѫ��A�=�6�����mmR��u��pq�T�1�m�L[@ Ջ���6� uMoS/[���6�+�P���{2�j�z.4/5Pm� 8sZ�v�v�$۶ܒ$��dv���UR�!r!�V�U�k��"Ľ����Z[�s�� ��5q۶̯|[_� ��]���rl���[U+�m!:t%�*�l�ssʎy��^f�1��jَ�@�Q��Z��z�����E��ej�'U����7f�ed�ҭ[�2L�(
����+ �-ù��m��k��0��m��=��8*�S_�Wo���l���6kj���UyUh�`�)�nŝ�h�4j@���*�U]ûv0ò9ݎj*ڀΎx��r��N�j��6�\�l5P��
�("x��N�FbZN
(ݑa�6��J�Ӭ��ltV�"�������`�	�A�?�l+��mR��]�(c��4,9շVpA��vϴ�l-��m�ٻ"M.���ɍ�YVMi�nv춦��JU]\+Z%������M�- m� m.���NY,����I76ڷ`�j��:6��Uj���S<�rgiU��	��ummͶ�I j��ImlI�Ŵ �� Hm�L�! 8�
�/VƠj۪�v�=�[t�����;�sU*��uu*��˭�ͫ.�� �ݪ@j^1KUuU*��)X@$l�ٖh��6�l�� m l 	���ė�����`WU-r��E�A�D��i����Z�\�z� �֛I��9��&���U �G)��W��� [F��n�.��R�V���k8�
�i���B�[#cժλ    �ŷko/F�UR��2�RJ�m�ƲU$�m�h��%��m�s�gE�@UT*+�6ڑ0�mmm*�9��=T�ST˻q��kv�Y-5@e=0^������ES(�<�Rt��E��6�-�6��iBq� {n2lf��)!�p[m��z�6��ua�t��=UUM��Ac��B��b��s+��Lh�`̇ij�Z*���W��t�ҭQ�5I�E�iK���90f�'2��U�*�ɤj몮�2-Epq��Uv���YKh$s���ڢE��(���_3�]U@m��.ڶ�m��v����`��[d"Z�Sb�k� ٔ�]r�T��`9�W�U�
��D�9X���e^�j��V.+��#�Z����wl�ln�,��l�gK)m -�[\�&�3ڤKv�t���GZ�I��[�6yJ t�N��e�m	7[uv�ev�vڪU�jC;��ul�T�N��kԶ�$���ϧ����Ϋ��h�EZ�l�J�-�5;�v{p��LC����5�[OT  Z���Rz]=�2PU�  bB&p���x�����U�U���Kb`B��ٛm����-��`��u�����6p�i�`�n�.�R��)��d6e���ӯ����K+��nQ��P8��
�˲�j�y6g�o�7Z�:G3�[@ �	m�/u����F�l�4�K[J���U�+�2��� *�p��]m�`  m�p3m֋o$�����L�P��
WK�eY��U!5T�t;3�m��e�,6ݸ��gB<�UUR��M���յU++�ԅ-��r��m�U�j MӢə�� ���nk#���\�U(��v%km��b{)��P1K��ER���ej�uʳ����
�vfs/5Use:1�Ij�vT	Vڭ��f����%�v��Uw�����C��T��RWJc���મc ��R����*ni҃m���Aam���PUN�%^�ƢYw����eZ�e�WB��YX\�"fv��A��J�Y!п���Զ���V�9̦D���f���i� ��Zr�t���U��vvn��0T��`�nrh��6Cj��Jt�uU�T����^Ѻ��&�c�xVy���;��tp6����R����N�� k\�8�һl�����N8,�qs�{��/�6���=��w��D����@���B���U?��O����?��6���R��� �h��?�:�Pڇ� �6���qA8/��$�J8)�t�@�z
�+ڇ���Ev����C��iw6���|P�CB	҈$���$OP:A�8>��#�v/��!�(X(&	�!�Uܴ�v��P&�� �@� h"��}UN/j�2�ɴ0�:�!�$��AqD�Q ����\R;LAz]�LBM1TlW��������	�T<TS4";B�J &	�D�C�@Nx*{*'@�����!�� �8�����d!h�% �-"�+� ��$"��;P`v�=��t(x = ț�� ���/������X2�p^�8��`&�У���#�؂�x.�{�!1�'��x�t��<8��|q^�����
xo��T҄!����m@�����	�OBC�;H,,�
��
�4��#�FÀ� &" IҦ�����v���qO !
'�/����r**�����u��������
?��A?�$P��I@���
�I��UI*�C��rԸ�ar[��l���M&�m�,�  $   UF��1[<�ܕO	6�4���(� ��R�Ǩ�:�$p�7[6����9f�m�C����Mtt�:{�ѱZƶ�>4�Vk�,���Zl�ki�m��h�      �`6�R�� sm�[@-�6�  6�ݶ����� �l�6m:� Xm�[4���$
�-�M�),��h6�i  ���mkb������2O#����[�HӝN���q�Q�ڻ	�^zY:����(�r�7�艥��O�&�yg��'�+�z��,��v�z�ys�]n5GK���f{v-r=JQd�m̅Z�n��c	&xCn�f�]���v7cmnv�X�����Z�.=��w�l�%�$ �!̫U=]h�t"��^�d��]�ư��l��([c� &˗P)�8�=����ӻ	e�s������"d�E^z;K�$���q��K���%�&LPc�omֻ{]�3�I�]=�5��
�P�*��ㇵd8el�v�� 9�`^Xd��#��r�_fI�2[d�;m��OC�E麈y����quoZ�^태�I��ku�L�B��+�g��4[�y`$��cc�)dN\�����3�xԞ̽Cڶktb�r\�1�J�{z�]]��2'*iz6��������� k� 3���SԥgH;�� r�up5� ř��ۀݎ-=��
l-� R��n�9���F��];[l*�˵�V2�f�ǧK�RP��zq6��s�����^�kb؞5�#iy����tZ0�����m�ll*�ҳ�쨑g��q(]�H�.�"vk)�22��x��fTkR;Kj�낊�ns��i�t7��^眸I�X���tg�����m���q'�&ŭ�z�N2�\k\�#j�b��6������$�r=ҥd�b`R�f��@�6[�d?�6�i�EN����N���M���'��t"��z�B
l �
b��$�T���a6)	.��˹#fM�ݸ��t��z�u�N
��X+��Y���Ɵ]u,N��ʼ���3�NMN�q	n�m�:H�Y��e�Ќ�g��M���gd�+;\��z�2��;v׮A,ls:�Y�r�;z�=��9��;�N��fT�q��3,��\6�=���=��� ���h�G=��a���֛��Pՠ�s9�d,9' �њ�]�9����;/g
�M����l��\9�����a�����ū�Wwn�7�w*��X�����{q`�۶�U�;�w,��,wf�7ۋ ��ŀ{��X�`��^��$v����ŀn���=�n,wf�wZ�c�)w"-D���� �}��{�x7ۋ �׺��+���"�=�n,^������7wq`��p$���%ݻr9���%�ո4�I�.�v�	�rv���K�ڻڠ9m˸Gq`�v�o���� �}��v׵��d�܅ܼ�|��14"G`��^W�߼9W���,^���zX[�nK�-ˑ`����{&�L�������Ҡ��^��$�d��ŀ�`�v�o���� =�mݚ���۹d#�`�v�o���� =�l�����=��5����m�C�7<p��
�ѳ��i�1�ޱɲ��v���v.y��=Tv��/ ��q`������^����.ǰR�D]�\%ŀn���w�0{�x7ۋ �7u4�W��ӗ {�ـk��õU�ڪڪT����7��ŀ����6�M&��J��H�f�W ���p�������w$-�#��]��9��X�e* ��ɠ<��E k$n��L�w�r�WaxwD�����l��<�\s�]��Ӭ�
��9�l�d8�l��MMw��ۻJ�=��h?��@^{)Px|Q�4I.Y"�v�, �}� ����o���ŀݶ��VD���YrL��dP��TjfN�n�* �f���U���rK���x7w���ʯ<���N�G��1�Es�UBT�SUS��L�ݼ�r�D]�\%ŀs۸������� ��~wͷ��۞^��eE��1�/�k�8pzϳ�F+s� ;���S�t%��s��� =�l�7ޚ`��X�w s�4�܎��r��7ޚ`��X=�ŀ��`�-�$�ܹ�.�7w�{q`��=��zX[�nK��-�rH�{�L ��� �4�9���|=��ZnK�Wj܆ {�ـ|�*U߷>8~�����߷*�R(AfA#��ow������C��"�fZ�c��g�2�jv�㪪�@Uy
��e�n�WR��<�+Z
-����D�@f�te�H�"v_(�;x�P��N���X�r��v1�[�ӯP�꨺c��ks��s׻F�&�8��$ˌ�����F�.�v�]lj�Z�ݖo<�hc����q;v�:g9宍��SjdC�g���]w X0������m�=�ۜO' 7 ���J�I%vF<�qH��@Wq���j��$^e�{�東��mҿƟ����u<�bE��$�K!��{�7ۋ �}4�w�0��{V�Iv����\�&w3�:P{6h�Nٙ29	rD�Ȯ��=�M0�������ŀy����7i�Q�$0�������ŀ{��`{��bnG܃w&��� ����=�M0����7m�c�Mܻ���C�g���Ѯ��	;�(�0V� � �w9�w&]��Rt�m�m���I3�f���� {�ـs}4�;�Kz������Z��U�~o۝�b�`�8�0`��|As`�o~{�U�~{ŀswq`��l��r\��V�0�����ŀswq`輦��wf�[w�j�ɀs}��n�,��� =�l�;�ަ�b*���iܸ���T�L�Y�,��z��J�o������r,W/1��ny{u���v����'��{�}��b�Yj�j�KqHK� �}4�=�����ŀswq`f��MEq�%�c��~ן%T�;��,�}�,��� ;�v&�&�pm�-܏ �}��n�,>T�)QL�(d�2mO^͚(ln= g�f)���ܖIw#���ŀs��`��^��q`^�Nޫr\v��r;���i�{��x;�ŀswq`�y���R��1�m�gsi5�۝�ѕ.�\U�]����ڊNŊ�Jf.W�z=�@_��T�e-en{'J �����v�r�+q�w��q`��X;��_������؊�vH�r\X7w��i�{��x;��ݼ�r$��"��ʕ>�s� �u��ʺ���r�
�H�,J� 
�K��]��,���hj'�H`��^��i�swq`輦�_��ƭ�.�V5r��@�Wvy��t�7ni&;�s��ݎ��&�y�"��pWH�rKw#�9�M0n�,��� �������i4�]�6Zv�8n�,���l�|`��<��� ���v�[��廑�Ȱw�Lϻ��s��`�n, �n�djܗ.8��r̓�{v(����{)PjI?��Ӏ"��V+.�e۴Zk�g|���n,��� ����� Ի,�`-f�ի\�,������{I�K�=8 N�[mu�&�dɱN��,�0��i):�Su&y��s���fVK�;Y:�l�Ҧ��q۵�u3�B=���Wb� 7)��^^y�ňyx�;��(f�v�z�ͺU��س�ᛍc=v^̝�֠�4u�q؉�d]�����{ڝ��R��?�tb�;V����$�Y܇n��!u�N���wx�ww�w���t��i�}tKD�v�!���l�8ϸ�kHݤ������ir���e�k��]h�Tt��W ����=}�\;� ��Y �.I�"�K� �}4�ʤٯ�}x}�� ��q`f����j;�e�������=8J��M���k� ;ݻ��&�仹r�>J�}�q`�~ŀs��`}ݼ ���$�n� �;�`�n,ꤗ}���5�� �}���F���Kp.�atGp ��=M'v��q�\t]F�Ʀ7r4�t)qu��.V�v�i&�&�g|���ݾ����;��X��6Ii�.\q]��0�;׾�;A
	B ���eFBd�"V	H��!�	J���ߞ���n,��� ׺����c�wn��9�n,��ŀs��`�����5{V��r������9ݚ`{�u�{�n.n��B�.K��)	q,��q{�u�y��]�lK����i��R�Ad&�oF5���`��_.��N6�vܙ�z���&�����pwRI��{���n���b\��r�ݻ��&�jX仒��۹�~=6:��l�{��s��+��Ji6�Zd��.L^�~�s���K��*k���(R�=�����^f��+�7�ã'|xGM�8�Q59�.�����;�f�@%�	��9x�I�U�E��pQ�s�3�;��"5��A���69:<"�4!��u·zyS�ζc��\:��F�3����d�5��n�쎜�;̰��'��H��^�CН9ǔ���b`�m4����CBB�f�,�Qц�Ӡ��ޱ.���`·LN9��ę�p��vt�	���֎��P���oF6��:����`�.(pW��6.�]���,��>PL��:D�/�x�Pc��Oz�=�)JR}�}��R��{b��K��-ܗw"ʤH)w���Cԥ)���┥'�����)W�߱eR
�
��Oݬw.89l�s��)O|��g�)<��~��)Jy��p┥'^g����R���w���;h	�g
��!��ۮ�c��Je�[K<OB���5�11q(�p×\h��Ӗ>y)JO;�߸=JR�}��8�)Iי��i?7r�������)JO~�3�l�j�kn�{��JS�����):�>��R���k߳�R��w�ple̙	�fY��D�$L�;�ʙ&%R��'~��hz��=�^��R���}��ԥ)���ÊR��y{��a���H<��U©R�^��R
^w�pz��;�߸qJC�� �ŀ�,@���FAaee& zX�E�@��r{�s��=JSH��]�����;M۹�H*�R�w~��)@HO�{��z�>���߾�G�~��v�4.�ʆǘ�E���ZOv�I�4<7v�]ۍ�L�Z�Z�-0:ַ��R���~��)JN�Ͻ�Cԥ)�}��E%�JO|����)O��?8Kn9wr;�U �AK�{���JS�>��R���}��ԥ*��Ҧd�}�O�m<B��b^Gp�s��)O|��qJR�����R����Ҧd�_�sa5������|��˄�ɕH*�R�w~�\*�U}��8�)Iי��hz��=���*�/n�v�W�E]����p�AT�����2��!���Л�2��)_�Bd������)O5|��a�N0X(D�,A���¿u�[R���7b�7LdP��^��{I7q:��	��� `��a�յQ,�E�r�j�{\$�d�Nn��c*dx�����(�ӫ��=���Ṻ]-��Rv����򬦶mq�R9��N^v��;=+k�8/ q�Ŝ�W�g5=���=q�͞�t�<�l\��H�x�gr�������y�a��g\��.Z�%��=b����e�E��;~�Z��V�1�?S�.��;9!1��n�j���!i@ڵ5�۶��y���6�Y�z1λ*��3[=R�������R���}�)JRy�����R��Ͼ��)JO<����9�����U©R���U �)<��~��)Jy��p┥'������U �F����6�R�"���ʤ��w��pz��<��qJR����~��)@���p┥'~��|o5���f���j���R���}�)JRy�}���)O<��R�����ԥ)��> �9,p�w#w"ʤH){��~��)@E�}����R��������3/{v�3 f@ˑ����Jy�y5X�=j�)�]����AWf��cZ}�S4�G]��BɆc�YvK��32�t�AT{���8�)I�{��JSϽ���d���l&��2��x"NK�D�՛��)JO;�߸=D��L��s"(�(Hg$`LDŃ��C�5)����┥'���hz��=��qOʎb��;z!Ө�CD�J���Mc2e�߸qJR����~��)Jy��p┠R�~߱W
�K�|}xZwq�-8E$�l┿��$�����R�����ÊR��w��pz��<�߸qJR�����wv���.fE\*�U.��b�)JO;�߸=JR����8�)I�~��R
��>��$��j�%ݻ�խ�� ����=��Dv��ጯR�8���t�܉�mF;��.,�AT�������U��{�)JRy����z��;�߸eR
�������HF����\�\))O|����'�~���R�^��T́�/}����d��t����r��nH��R
^��>p�D�{�)N�8 �0G�M��<���k�3/��J��3 e���M����&%Ը���5��93!2�oZ�d
R{��pz��=�߸qJ�6I�g��3 f\��r%�q�)���T�)I�{��JS�=���)<��w�=JR����8�)I�~�Y��hY��B�۵�7&��kEl�]dP��0:ݷP���g�e8�yr�t���)J{��┥'������JS�����)<��~��)Jw���9�ַ��R�RK�ʤH){�l�U©R���ÊR��y��pz��=�߸qO�� e�wrw�����re�&�Mc2O?}���):��~��)J{�p�T����>p�AT�߮��&��n֭�g�):��~��)J{�p┥'������JQ�'b�ϳAT���n��ܒ&�#r�R���{�)JRy߾��z��>��T́�+���k�3#p݂I@C��Wazm�.��{v�ݻ<�\8�b+���!�<	�k:K��4�4F�֫a()<��w�=JR����8�)I�~���JS�=���)=;3�m���֭�xo"���z��;�߸p��NJR}�߿pz��>���8�)I��N��e�328̹�^�K˻�����┥'�}���JS�=����I����z��<���R��^�~�i��"��vJrLU©R�o�qJR����Cԥ)���ÊP��Hq��{�5����N�P��r&$�&��kg�);��w�=JP�O�����)JO����R���{�)JR5IR�����SA��Er���r三v���P���3&]�M\� �����˲��AɰÆs�i�5u���m��m\�w<5�Z	[˗�]k�y�ܬH��Iz�J�G�,�1û�Xvq�B��<j��]��\�
)��H���5�u�����a"L�L;Z�mVy덪�`���z�헖�r{�<qV����s�n�yǷnD�vtuݯ;���#	��n{�{��z�9^��aȵsZܯ+�k����g��fi3��m�m>�4^���1!Y��{����>�R����)JR{߿}��R���~��)JN��︽JSH���mKq�d.�qeR
��w�=JR����8�)I��}��Jiw��U �AK�}��$�&�܅�v��R���{�)JRw��}��C��d����ÊR��}����)O���%����,�AT��~��z��;�߸qJR��}��R���߱eR
��y?^���%ƮX���ԥ)���ÊR����pz��=�߸qJR�����/R��߹��|f��um�cÜS��Ծ���	�ۍo��e�룇�#��h��i
��m���=��ԥ)��ÊR��}��qz��;�߸qJR����Z�}�sF�V�޷��R���~��0O�B�b`b�JB�B!ࣷ�����?qz��;���g�)=��~�\*�U.��֞�e�q��˸����}��qz��;�^��R�������sz�X́�noR�d�_�f�nݹ.FJ��&Up�AT����*�U�{�pz��=�߸qJR��~��/
�H߾.Ϣm;r�je��QI�{��JS�=���):��~��́�}���́�+�vIC�<J�r.��<��<���ZlD��8�b28Ɉ������Jj�k0#|�}o{��{�p┥'^���^�)N�׿g����߱W
�K���,V�rۍ�z޳7��R���߽���~ ��O?k���)JO~����)O|��F��_/'�����c�W,Eɕ\*�U.��~�)JRy�}��CGc�x!����S]}���)=��߸�JR�g��"21�R)n�<�AU��T�[�����R��߿p┥'~���^�(\�K�;�L��2���:��3�w�M[��=JR����8�)G�A�8��~�q|��=�k��8�)I�}��J��}���-,�k R���ι{v��לp��.
�v��lr7��v{.��������>�Ǐ��\����&&"U3 f@�����c2e����┥'�����)O}��R�AK�>ߔ.�r\�� ܙU©R���RK�	8́�vwRk�3-��T�Br�=��~��'�a�K�Z���b�ywxR<C��3 f@�;;�5��ٌ�߸qJ+�}��qz��<��~�U �AK���.K�;��`ܘ��%~%~���R�����~��)Jw�{���	�F���IR�!�I'K��P2����&��2���8�0f�ݭoy���)JR{�����R��I/GoE3 f@�;;�5���{6�3 �AK��i��L�%��,-آv۷9�ݹ=��[`�ua23k[���1�y���s�\}?�V�Y�Ʒ����{��<��~��)<�Ͼ��)J{�p�~�rR��}ަk�3.|ׂ9��
$����fT�'_y����(������)>�߿qz��;Ͻ�\R�)JN���k5���֍�o{��)J{�p┥'�y��^�)N��~��):�Ͼ�\*�U.��֞�v���%˸��?�L��}���JS����qJR�����R��	O���G�)<����չ.Ic$�*�U �]}��R
J?���������R�������)=�߾��)Ja��G�K��TY��A�k�6\գ1s��pu�ؙ�ĝ��m����#k����UP.P�ëc��͑�(���tb�$V!p���q-oh�\���:����tu���F�I�D�gC��9Ɩ_�����z����F�O�t�4��e���3I����E���r���w�HN�NZk*R|�U.չ� t��5k)�kZ�)���M7\����p�7F����kfٹ8˖#�12�S�[S(�j�ʼ�in��0�fP�y�ha��a��üָٿ9���R��$v.�b�������/[2��j�jB{�WjD�Q�]b�;yTD����iM�<�s��u�@�z���gX�0qS!E�/L\L0�s}#�5��F�G�l����֎p���[�zqu��H��.�xwl�,��2�]p��-\��Kh<�Y\U���P"vp�1p7ͦ�0�`��d؛*���	��ː��;���I�z�G��6؝   H @ K������qj�`�b�QА��p�m���p`�*֘�ck*X���u���[�[(<�;awg�H-@mѽk'\=��ʣo��Pd8i�         -6(�g : :��   ��m�<m�  ph� 8[��HY@vq��}�Ãm�mm�)"�;]0��,� �q!  ��PPM�ͨ��8l�HΚ��oNw��9F�8b�^�$n{Q+��kp��{M[�8Ś��(It7s��l��^�j�umѶ�GK�^��H8��ם���*�J��7�V��I\ݻU�^XM�jx����p;y{:��v�"`�Wb�5�ݸ�w�1=�;cî�������Ř�l���<0����[m�n�Z ���S�Ѹ� j,G�i@f����`�W;��)-<�1�*�m9�:��Ojd6�z�<��ŔZ5�t����9�m��n@�m))`��\�6s���m姴���3�"m֒���X��}]Tua^l)K��]h�PZ'��}lk���!��+pzݷ#�w[�r૪��".�㭈�y��ŘQ"�$ѹ��!�S���m�q�k�sf��I�����0V���Ŵ��W��r�n�0ueV��<��g;�i��v����@�N�I�'@��OBm��K�[aGg���i\���kCH�D.����(ƇZ�sm3���vS<�l������@���Q��GQ��2ݟ�o�p�A���N@b�zy��F�q�-�;	X�k��#Qu�@66�����
�
�v��p'C�''=q�&�h��x�XN3$�ô�h1�'�RvU������Ju��l^k��62��2m�qv�6������p�
+8��'d���(]΍e;'9;T�dL�]�c��H�iz��	�[I0�$tI��"�v��+��[T�T�@��Ђ�U�q]�x�*'� �*lE �	�&�@^Рbt  gm�-j��n��ky��v�$�q�l�9_nju4ēN��U�ݭ$�H
ڡ��[Oes�K�N�����ڝ�e�OFln1�m���켣���k�����U�`3#��O��fE�D��.�Z���I���2��
<d�v�g�l���v2ar+�|l\���\��5�qc3�uc6��)O`�k��\$3R��c+��!םN�Ӯ�ؖ�u��;�G�T�RT��^��N{=S�8�Lv�\����ѥ�ꕭ�nv۝�`s�up��9W=����':�y�J~JR������R������)JR{�n�nf>�3/?wE3 f@��7z%�.Ew.)%�rb�H*��όT�*��JR{�߿qz��<�߿k�R�����b�H*�����c��rܻ�U�'����^�)N����?,����I�f@̷vx�d�j�?�U(T���&��f@��Be���)JO?}���JS�}���?8�s{���d˟9������L�x5��R�����pz��?����qJR��~���ԥ)�}��┥']���y��-4v�!���l��q���]:�b�E[&{��ػ%_?~���Ҝs�v��vo{�Cܥ)��o��)JO{�︽J2��v)�2_nn�k7��	�"#�-��rC �o�qrR��"�E5GY�:����a����H�	i�ܑ��;���n���:W�2?C����LN��I�v���7�_ ��۱�2N��<P��`7G����QK�2�ܒv�}`n��@gٻj�M̒:3�(��藘��12D݃o0	���7�&V/�.ٻ36ߟ��q�󬳄�P6|�hm��SIݳ�t�:��Ӧ�n6u�zqu����ᾍ��[.�M[I����_�\�vg�~o8~���j����PB��I��Ұ5���������;vx�3�+ ��hQ�ڦ�݉5�;7g]U����f����=���D�2 ��Ϲ������~��A��t�>�!DD����~L���v��7��j����PZI��ڠ3��	�v&��I�m����~��T^�p����&� ��۹J��Tպn�q��G�����O.���pd@M�˱=��N�5�gJ�1�Ҷ&�'��K�vn��72t������߭X���C�&TA��L���m�ɹ�v��@o��Հo�f�������13)��b]�fn����ϳv՟�����=۽v��k����u11Ps2C%�����W��?o��@}��v&_&y�I��f8�02J�T�!!),(`�%2�dA�����/�ȯ� ��H��`^[�OˋՎS�6�0��l���t��#?w~��z}���7�"%uE;���j�%E[��ognzݎ}�9�����=
�og[sɛ�{e\�*\�4�:NĚ���0	�p�ݜ��\�����;s�9҆�O�&fn��d�Ip;��������>�ͻT��	;I�&�l�ݜ�/� �ݙ�Ok� ��R�L4���2�E���2vI~d2_�{�P�����(.HI?�����.:T:�w�wO1@{�ݻ%�	vmq@{�=�`k�6(���L*C$�bA*�2���G����[�Y�ݼ�a�#�Ӟ�ac0��\���u� *6��V�n�)���
��Ik�n�M5�:��Xڶ��c�1-��x �Ϣ��U�Z�0�VE㛘1�.�C�nu��t���t�����w����L^�;vS���Y�8x�8�t`X�m�!�3�6Ƥ���cg��G)l�����_>s+�d�F�m��󰩢hެ�Gi�{t��fu�--�
.�ʋ%�.Q�m��t���`�y�m/3u��ܝ�R�.��I��M��,m=�?�����e����$��&�&BJs~�S����0L'S0�1%��9�c2\�BHfs�7���gu��(X��;�!@��2�⪞���lP��n���L��2BP����8�����_��%r�6��Iآb��.fL$���vf��l����7f������~�4Bx�0�3���p�9/ ������� ����{eݚ�e	Lm������$�xٺY�۶��(Z.�$��YI~P�)P����O'b��bi���|���	�p���m2nd&�ݞ(�NP��%LC���3��:��5����<�qS��I�ɫۻs'J���{��$�%�!4������u�;̻����7{�]���ҏ̝%���G���������n��V5m�N��M�=�=��o�5�?2Hd�2n���`b~�8~b&���L<�I@}�װ?2L3/ɐ��Ͽ��I���`���3e��:,���U�֬�)�]��e�趫a��r�؍��iۮYe4���0T�ucj�9��'�Ǡ=�ݻ}��3s0������>k��f"T(���zٛ��$��1H��?�o�����	���WV+���O���}���l�o�2J�M	.fd%GTo=���`fc�'���!�&d������&a&��ߧ��?lw�=��v�$�ٵ��a�����y�2�sO`o�5�3~a�n�W�}��p�r^���lbi��'*+���.�zw@���9km��]�ob�	�f����$���,9q�n�˃R�<~�}���p�r^<�_ �(�N<��Q�]�&��N���a/�fHa%��~{��~zٛ��3�%��!%'�Ç�"`�N��b&bJ;������|��3 ��+�_���,�.�UO`$˄�$%�;�@fn�몾���r��ZX���p�Q�I��(Ƚ��J	Hf�>�y��6�����R�t�;V��{vf=�=��O-��=��.;��Vփ�wm�c̛��l����p�y3G��KI��њ:����\�Z�-g[�U�M]�΁����3��x��|�M�22�fp���7u��DK��6�ն���e��~�v}�}|}���7�:W$$�$�d�$��?(�IrbA<L��S��;���ٷg�ffw��w�O��ĨD�Ҵ���I7�M�! d�>{7����‿�6Հ̹�d���>Ӻ:&aǙ�yQ*%�O0	�p�ٳ+ �[/�{�٘i%�R��j�>�}L/�p$��)���1�������>�pUUR�\��L<9}u�Q,�<���ڐ�R�fM�YJ݅�.z6(z�D	5��_@��e�s�i�6�����Dxzs�Z��T�<��s�'j�׶W��I�C^h�w�#�Ѯ�E᫞��O'gMf^sm֤�f!���w�����2L��k��H�k 5��k�C��WaxwF��\�ݰ�'�p�U�cY�2n��Cv�n���;���fhQv8[0L'��������~��Ձ<�_ �}�0	�p��K�q�*C�<˼DҰ7њ��fd�̿	�77�]��z����I.I	���x"!��6�@��n��gـOk� �͙X��|{�+��G�J���`&I3�_�	����P���Ձ��נ�ɄߘJ77�]�����DK���30�,�ٳ+ �[/�{�٘��p�~�?�E>�0�Z�s���\�8��Y���m�L%�OZ�K��c����ER�Ê�*@i[����|������w�3 ����2�ޕlt$���;)$�{�=����>|�iMjM)�T�2Zɖ32�!0�����P�޵`nFk�!2a�'��q�D�䧗����z�nm�?&fg~��z}���;W��YBiڡ�M�I�
��&d�{��X�����m�~d�?gW-�z��
	�<˼DҰ7#5�� 3g�z�������V�~�??8z�XIۖ0���zl6�ݸ�p�� y�mn�����������K��gf�{=��`o�t�/�ʹ� 	7�tS��n��Պ�t~�whn�y�OG
e�I��v���7����ͻ3a�X��[m�ڻL�ٳ+ ��_Kð�-e$�Jz�(ѣ�h��6l�\�X�^��So#Q-e�4tl��������&���މ�4�R����f�&�n��E�o�ÁA(t�6��t����9�ֻy��v��04Fk�L4���4Q�x��:|�v�����u��q��Ogo �m���sG�Be4^��vf}�r���W;Orͦ1�Ȏ�#�La㛶e��[�z��n���#-NIA�:>P۽���΍8�K�\7{��(�Ӆ�Z�.�({Xv���y��XQ�$Jr�����F�H�ָ�aeE���s:=5����(CNQ����F*z���4{���Ӳy��u�l���H
JJX)8^re$JN��	S�F�qLc{�L�~�lkCwtw'{�p��,���ɡ� HC&��N��ѭ��q�#��:h		+@a�y�kiy����+H?*S��`��"��6���X ���`���@v��HC �.k��˰=�<P�5C�D�;ˊ"e�fՇ�2d�۽4{7��ݍנ_�'�ݽj�3yp�$�"w&]��5�=�l�E%��ٕ�H����~F�ۑ�����\<����n��J9���8�e�� V�ɗl~����~�L�-2�^f&��;����6Հn���ɒ��g�ـm_�ş�P������;�ٳ+ $��w�3 �I|������R*ۻI�I �}�0	��2n̬\����@�lT�\L�.B}��]����{���/2�iRb*�v�#9�Ł�j$,0�l�؇5����wڕՊ����Cv��H��
�ݽԾ�����fm����?n��	`� �E����۷<玹�p�ݮ
�v���wI�p��φ�$+_]��|2�JXӛg ��ﲰ	rE�7۳0	#� �i)\�I�.�X�co+ �$\��wwf`G��2��ʅ��բ�"\O1@{�ͻwgJ9:O�wu���� �I�&Չ�nմ6�y�I��wmX��ǽ��`|�5��N�;��;���3�L�\�p{w���*��C�'9��{�_~�?<�����v���3��P�{�:cv�v�㪪�p#��T�d]��@��u�ւ�['d���i�����юsMN����6N1��Ɉ��F�jy��a���gj�p�,P�r:�Lv���xy�{x7Wa�����RI����w:�=���{f�����Yf�ZlMn��>%{\���nrui8m��}���ۮ��:�������nPn��������3��V��hw]����]۷;cK�,��㬐nZ�B�	qYk�R�Hc.�ɖ�R*۱���^�����3 �8�����V?s��fa��0D�P�3n�̄�wt�@}��j���دə�0�&BP�~���H	�ȉ�&&�����p����%� �n��7v�r���!��&	�fJ��O�n�������fm��:P�5C��w�x����V��� &\�&�7z�����ݙX�j�C�o𩶝"��Y{u�Ó���Ѧ������kv۔�݌ۭ;gr��b质��evU�� �n��$�=�3��ՀK�.�K�j�n��;��������4�,!0ى.&��3-f^d�C$���޵`c�tP�ͻ�fI�39����1#�u1*]�$�>�޵`k��Q̝��޻���|c��P
y����a�̔&K���͟f��`s���`{��%r�7$�1@^{6�I	.�(�7�\�p�1����j�i��	m�#���7=�����[mL���P��e����*Ֆ�bO0	#� �ݙX�"���a�'ـI/�|��ݵn�g ��̬\�p�l�H�ϊNf���B�P;�
"^ffՀwwMy��d��~fV��I��wO{�֬�ʅ�+���vX�|�?_d�f��?���X$��{jh�wc�Q0�����wgJ�N̾���}�πwwf`e�8�ۻhI$�~b������d����w6uh�F�<��=t��R��M;T�t��g ͛2�I �{6��|�����t�P��$!����I ��f`�Àf͙Y̝�~8��~P2@�!334no]��8lٕ��>;5+��)AO<LI7a�ϻ����u� �����LQ �x�"�!�o=ٸ�\Vrĝ���t��8l�*��;�l�޻3gJ�n�A>zK�$&�o\�O;dn�@z�{^;v]۲��	;��5�k�盜\��W�}m��wf��fm��:rJ�>�޵`o.V�r�N1�r`�o���O�����wvk�L���D���?L��0���y�?�f͙X$��{}�0�컟�4�S���;�����U�}>�`�}���l�H��%n�H���"�0Lm�V I#�~��fϳ�wt�@^nm�Y���
 sfHwYmD9#+;i���<<�yZ8���[����s�Ul�\����	ei���IkDƳb�ӷC��]�؜��b��a3��u�v8��.uu�M����[s�ͮ�m�-tcp��]�s(��6�c���;c��x��d�t0�Mκ��ѥg;��c���`q����g;T#�cػ)��gf`[�v��w�k|��t̗~��ݏ��)ݺ4�X�W�t�{;s��s�q9����CY:���vI!�جu`�m�����}3 ��Ҁ���_�%���4{�`h�PU�-4Ğ`G�6e`�:��۾I'�sw_��P��<�1���w��X$��n�f`G~�T>�Q*����ڰ�&L���@�1�~�4n��v�Δ�d���� 4�W��+�I�*�V$� ��&`�d�wuq`{��j���ؠ=����6ӕK�\��ڟK�+���r�v�vwa�K���κ�nfn���Ҁ��ݵ`k��rIX�Æf��`���߭4�[�n۾��2�Ч� Hxb�)
�� !�WW���{ޓ0	�e�	]֮K�
T�m1.�LҰ5����۳�$��d�����=���~,;�jp���!<L��{v���z�sbÙ'fHd����;1�t��<��K�7`M[/�w�lX�H���3 &֨�l���P��m�S��s���fh{\��ێ��K��/���~�������}rFVEۤ�n�yo�,\�p��f"����.X��"�%i;�o� �$��Ifw=������۱`zT.�]�m�uJ��\����H��K��q32��	�L�2��M��S2fJ��C$Udoz,~�>��(��h-�����E%���K�%�������{��߭4�UiӼ���}݋�2Cˣ�������	#� �˗��V���i_�:�k�v���.��1��a��ێ��sm�l�m}3��R�[�ӻ8�.H�{�3 �7_�ВHp��;�����P�'�ӵNۮ��L�$R_ �W�,n�*�B��ۯ�
9yr!�^H����_ �u�I9\=�3 ����V�wWrH�?D��4RA{����߿R�/�n݃�fm	$033$����C&eDV���_\��yQ0�3Q`n�Ҡ?2_���3~���_ �u�պ�lbi�e����/]f6W#�;�8=ny�y�v�{K��x:˵n�h��+�ۢ����I��K��� �NW ��n�CcAt��Nn�ݍפ��3��GoE���J��ޓ0^�W)��햝]�n�z�"�7wiP7&L?���`wGs��d��С@����SOa�2L���j�������z��3�3����x���̨���/2���۰?2I���=��Ł��J���f�k����N�Ir���
Kc��b\u��4Xlp�N6k�9$0xBbClБ�d1k#dd�ḧ́`i���EhÃȗ:���:�5j���P��Z(�F�����#@��wxq�ؾu�����l8�mX�-�������,��t�v���Ls��c$G:����gfu��6h�kn�A'az;6��Jxk@^6&e��Idd��}�	#��&��4��D�)���!tDm88�U�&a�'�A���w:l�']bt�p��;����<t��gÇ�A9���B#{:s�,��l�N�i�S�<!��+oLs1��A%���3�n'T�]��]��j�Y�8�ER�]�C�6���goZ4:QTɚz7�.��+8TIh��&)�s�o+��*ԕI��::�z�G p ��   �  ���;zHβu%�;6q5t��4�M�d��v劫���둖ݼ>81�hԌca�7Oi..�c+�s�Z�S��v[�닮�-�s�Z�@���        	� Ͷp%(N� �փE ���`  ���l�[@ À���� ��� Hp�lknA��Q���
Qi��K)J d$80`Z�a $�m��z�&6\�	j����������ݔe�����#�v�V7Q�y4�OUm݊�]n��IF4�fy��mt�-�v�sR�mm���x�6d�h�����\�@�r[�6�K��i�ϕ^� �E�G�\<�������6ʄNM�֓��]k�	;\�U�żd��f�\�ŽJ��L`�r�������s�)�)u�n�'`�p&v3��� ���U�s)��&+i|E+6���*�ʦ��6m��4u�9;��.���h����s�ۓkZ�����2X�n���/ML�Mvۦv6�U�$ە�X��ڙ��X�JێFJ�ºѺ0y�D=8��t�۹v�nrq�Zy�L	�m�������jq�ď`�=[I�#��60�[gAŁ�6�D$x�*Bk�g��Ǒ�u��6����p<vM�u��h�_Zz��8��y9�ê����G��\�<�Bv�*�W���gf���"�'��f�ٺ3�I���;rP�p.���.˦'��rv�]��s�ڞ.��:�ȗ75����)xi͸�7[C��qJn�M��W��,�5؁!�r�mv�n��Z���g�*v�R�l;n���]m[ax�V�U��6�`��R�����u�=�����a�{ ��(�\8��	^�81�VH�+ԷV�s�]���R��U��,�೎��=�.5�lf{(�{W���+��]`��!5�%��+l�Ӵ+�tdp�;t�,�]u.��ֲ͖��7� �@���1C�H8x &�E=�o����v��"i� 'i�Ҵ��]IRT�/jbhG��n�w{���U�籧��sE�n�z� &�p%���d�z��7n$
٤q�mttx�FB��.o]uv Ț5Ɔ4�*��usV��
]0ݦ�m���n�n&��+�L]���6��Nj�No^��:ɮڲ�-q�����]d}��p�j*�]�56��l<J����n-&�]��cfs�%�jE�C�ӌ=]�����YlD����l�c�{�ڣu�4���n�ɹ m�\	�`8{\����͎�3���<=�:����$[���wT��;�I��n�ү�d�{{�����
�<�<D�i�M�|���X�r�{�f"����$/�49�~_��T*"&b"m`���ܮ��3 �I|��̬ �H<��bA҄Lʠ��!~L���߾�?�������2�	$�pvt�t�?֝�i��$R_ ｳ+ �NW �와w��|U�	&�7E�h�n��.Sn {��K��J����"���C���(���w�n�yo�.�)���ݧJݷx�g�X�r�wd�E%���qۗ�J�n����o�U}��p��'��1��07"&ӧ4U!,�ݨF�h(K{փZ�6"v�/`~T�|�
��]���@}�fڰ5����-�V���u�3�&`)/�U����BBfٛ֬��T�Rjc�+j�o0	��;�l��$���3�&`ݸ*�+v�'C�I6����ZX�ɐ���{�����v�n�m�������̝`�W;�^r�X��k�$����LgVv{`ќ�x�g�3��.V�K8`G��3 �I|���~L�0Ç�'y�L�܈u�!�^���v��w;���fN�����=/mD�'@ۢ�i�"��~y�~έ�քdB�=N��N2���4jB6`) �L�R�#v�`'l�3d�	!�}ќ�۝�`y�t��& ��x�/2��&I��[�`wGs��n݇��d��!0�t�=��Z����J�n����/ �I|;�f��@}�Nk��?�k�'��	]���pk�g�D�n:�y'���a�nлR�7n�xT;�aj� ��[c�Ӿ�����0	#u����u�a����;����~HK�
��n�!���K���^"�z�{6���3~�	!��w?�R�j�t:t�m� ��?�� �I|����$R_ �[r�V�V�ZI����ː�a.��z=��`n���ZI,�J�~������m�m\�J����f`)/�gc�x�K���������6.܌�^F���ݞ{����B�mi|'�ȏ����b�]��D�T�(ES�>;��i��av�|������v9/ �O��{~� ��cO�.]���+q���}� O�� �)_�濟��O�� �I|ҍwr]��_�I[J���-��=�l�E��v9/ ���� �(��TDJ��̒C	�C&a'�f��Ѽ������NW �nB���+C�ؿ&�`�"��N�������۰!�Y�`�/0�8�P�b�t�k횴kzֵ��SEp-��;����]<���UT�6WeY��d�a�뮧38;;��n�N��m�ڠ�N�	�6+�FEy��(G�z��W�;s�Җ�s��T!�4G�N���r�9�������sʙ�r9ɮ������1���vc;���n�6.���3�����ܝ�n �YT�5l��^���V�i4�v�^ܜ�-�o,�l�Z���|P�C4 ��T�IAY�	
AD��� VQe�)A!D	B���nޭ[�݆aUD��Η�nyɵ�&���]�)v�����Y�,�s�pFV��i��~��w���}�J���Ϳə�����կ�By�LA1T��gJ��L���$$�L330���7�����/읗�=!wV��ۢ�&��;�l�^�\;���dp��À{�{j�%k���9_�(A�P�YP�c3b�����}�J��I�ٛ�X��t}M4+v�ӥbmp��C �?W�%Y�����tr�=���uT�ظo����b�І���S��6ݹ͈��ݹ�[c��k<��g�rc�թ�k���|�7?�HM]������{f`�b��y_��-T��	���u�=����T�"�<S���3	@�$2L2B��K����7��Ł����'��U�ӥht����y�K݋�u�����@�Q4��MH;�wR�3ٽvx�aRw�����)�I����`d�pw�3 �� ���ۖ���N�$�i�zNW )��L�!̄2�f�|>�EnV����t?�,B�y����ゝ���xn��p��kkn�FM��;�=� ��+	*MS��T�u�o�}��ظvo!ɛ���T��GD����y�S����W��k��H�4B�4�+5j=��������6�?�ݍS.<1*���=��i`o�iQ̗�$2r�p�.�!#4 zu�%R)Vb��.������^�~�(���_6UB��"a�⨰��~��T{�����ؠ�fI�ݷŁώ��̢%L��U�6���&C&d$�!�{���7��,{���a6܃��wmF�0��v����1�r��[��pp3K�v��n8�CCe�m��%���=ټ�='+�{�f`�]�J�ڴ�:ui&� �~߿g_�1C���
�P�P~�ߩP�������ر�� ��3T��v��6��C2@ɐ�f��z(�N���l.�J��:��I�\ݛ3 �� ����z�h�H1pV��U��%�8�������u��!�(�Zv��n�]�O0	{�p��H�1$�!0���������=ٳ0	�tN1[I$6ВI��F6���i=�pK��g����	��7m���pPxtݗI;Iұ6����'��p}�����ßw�����_zUB��"c7��3����s�,$�)���7?w�??w�=��k��s��+�Am�t��p����%���7�{/ ����'��U�ӥhht1�o0��$$�	���w���d�=��ݥ@d���7ƻ��۱$�S�I6�����:��"2?�"�}��vr�O�� �� �w�6�,������㴰��u�^{=�&�v����;�j��"U�+eݗj���[OdL�P��-Ԙ뮄�%/Ngn��v�,E���.��n�'�*�0 �ܘ\�)�(�@T�Rs[�N�И����{"��kp���s���.]��6����\�)m���]�˻vMo<=���ۛ���{x;s4�[��ڮ=Sf�+��nG�ծ�������a��w{�;��k�nu���	��p=.�;ez��B}����<�M2%-#^޹ Um�RI���_����p�٘�ظ��e��H]դ�5N��ӮU��{�]��BL��#����p�?�� ����7f�Q�Hv���	&�|͊=��{?&d��;�Pvw]���;��e�Q2��ș��� )�a�s�}�߳��{��A��f/v.=�۽���QC�[VMM=��ݥ@~fK����w���zr^�(��~v�ݶ[V��4&���n9�y�PjH�t�I�6X���W?=���w��n�UI"��U\���@����Xݝ�`k�lP�Nk�I2�ó��ٯ�'N�C��$�����_3b��I43ZL�ɞ��{sv�{�۱������d/���~٬��&
�ZI��&�^='+�d���%���;�-Ɔ�%m��r�?����bUI �}��vr�?���`�E�7�{/ ;�WV���;ʓN�Ol�^ȸ��e�d��6�_�����f��r��z�0�u>�����(]�n;mfR@,����MF�ĩ/ĊTRE*�*)R�̷|�;C�)ws:>�E�zs^��ݥ@^�6�?�݉M��&�[�bMp���&���=�v�n�$ɹ��0�L����_zUD ���&�����@^�6�ē����Q!v�������r���&vPFХ�,)3�Fq�1ü�:�{�X�.��u�cA;�3v`�8�`l�Ǧ�:��;�˭��KV��M������+F8��iIi6�]�<��1$���6Z��:��A���2����ìz2��9����١S�n���j4jÝ��.�sI�('2��H�gcA�&��A��' �;sA�v���B�Hb��tF���.h0]� u�͍��VSF�a�E��(�t8	�e�b`7K��lt9��u��-hBsI�#N�����D�\EL4�)�$&_U9�"�C��%�Ha;��#wFgg#k�S��;S@��mS�x8���1�D<J Jq�."(�H� ��T�+ z�� x�����g&�${/ ��{W)��+`���P�ͻ_7b�Ͻ9�`33s&f]>�+�}�����`�]��� ��E����[���Ԩ�f݁ɒ~�Y��l��e	}��+ڍn����m�ۮL�T�hчQ�Ү01ݶ{l�r���±1`o�w���ݥ@_�ʹ�ߓ�8}r|������:����Sv�{v�~d�����9�z(�Ӛ��>训$Ʃ���4�g}�0	{�p?W��&C$32��;�`vwR�=���)"�&�;m�/d\;��	�R��$��i3&f���\�W�=Y`k���3B��%C����{�3~�e`�f/�.�/n1�ݴ�	�У�	&��n.�i2��Vj�\���i&�m�8�� �Lŗ`№ɓ �w�\����%�E�2�6<^��\�Ct��cT$�{�٘~�U�%�E�2�6<n�W �6B�[h��X�o0n�o�f͟��2w�ޥ@}��v�lEm�[��Q;��x�J�)R_��G�;�M����*��۰5��bՏ�)�	�B�����s6���M�f��ϝ�@[���`;&��a�2w��n����a �Z嶅M��oZ3s���� �+Y�ܶL���X�n��.�,�u�-ۤ��A���7�:��q�FKm���:���`�x��
Vr�BDa؍� �Wd�Z<Sg�v+���9h�H�fmp��7GS����s�گ=�t{=��h<ǭ�0�5g�m�r� �l�����yhێ�6�v���F�N)^�N�ē�뉣=���}�����{���V�Y�q�TV՘헅޹��<�����vXx�x�p��`�}���w�_Y8I���t�����ـK�e�v?�߻a��r�Ϣ��hV���14��_۱\��|���;w�P}�۱�2��fsϚ��)�"�A*���>gs�&��p��3 �� �B�'+� +t������	�9\����%�E�dɸI'����`s뾧�(�P�L�͢Ӯ��f`~ظ_}#�;6r�m����1�sY��Ɇ��vl6�,�š�����hݞG����է���nx�D%(���n���lP�{vl�m/ɕ�&�2@�L��@fo~��~S�x��)�"&(��7���,IL�Ը����%�b��+m���'73U6�6���v�d�~C3&�a3����7�l�>�	� ����u�;�0	~ظo�#�'�r��j�B����t�i�/� ��_�tə~&�����|��Ԩ���`{��|5HI4���e�R���
]�rWfbv��쭸y|��u���KC�bMp�l� ��������������ws�x@Cʒf�����fҦK�̙�HfI�ٻ�`s��P��/oi\�Bh�4��+N�}�:꯳�~�/��	���HNbJ��f���ebIRdəc*�}���;s�P�7E	�Z�fl�n�{�]T(?�*�I��3z(�7�l�m*�fm���-:E4+�V��I�������;�٘�l\��Uo�_1�l.��r-\\�|�n��q��\�%�5Í���݃���٭l�h�� F VIR�i�+?rш47J�K��x���8wvf/� �["���@Z��M��I���3 �틀f��`���D��"��%(����'�;iX�4���cM����pղ,{\8wvf�ݻ��6�a�r"b��$�g�g{������=� �ʅ��CXCU�	�,m!`��&'��i�+�b�Ƶ/
$9*�Ck��4��4��h\�6��59�Ff�����L�g}��;Qf���LLÕS�uW�{��U ��a!@����)E)�<��s��g�~� �["��J��6!�@��aE��=ZM���q����ۉw��O(��|����v�v.�Un�[f�'ـK���3Vȿخ�}��p�����Wn����y�K���Q��-P��0	 J �&@��fI����g��ݙ����b����$Quwj��dXz0��I;���v�wE�XÛ�*ޭ�ѭk]o|�U?�� *�I&�mq@{wz�f�y���DU�I��U?�L��٘�l\=׿}����w�ʻvD�	�ǽ�Ǿ�8��jU��q;v�R��F�yX8*��`�����g��/�[��;��]�6�Y��;��e��yr==-g�S$�p�\v[[����-�]�������\�S�LY�x��G,"z�V��-���u:��e�g��=Qf�fqa�$!�mo9�(���6ܸ�g&�݋��5���]�FvI'Tc��l�ͶmGR��������&d�b�#+א`a���;n���O6��1�����j�kF�۵����HKUA_�y�ݫ�i����4�:�'ˀf��`���;��0�۸]�h�	�Ҵ�8^� ���ݙ�o�ÀwhD�����M_/�� ��\��}��)�@�)�����@y��~�_�J`yV�����~�}�l/vG�vk� �7b�]�hN��m���.U"� �! iiI�{��|����wwf`͌h�;]���Xi$���iz��G+ul���G��ӹ������;�.�m�m�}��~_X'�Àwwf`���=+H;�j���I��}�ڴ	"��*Gc�� t���hP("D�fBI$�o�����‷�ݛ �$
-ZM&���$��ݙ�Okҏɓ;����`vl�@{3v^G�yxwַlֳz���
��� V$�HL����(tw��`o�t�>�ͻ��w�m�:N�I3�f��`���;��0	�p��]]�&��gg�l�m��wn���۴0�x�S�c��i�6y�,��r�"���/�}���}��}���@�U�2 P)�d2e���,�����w�3
d�����wwf`uÀf��`�r��Wg�I���ڷM�T;o0�=��}��~M-�Iӆ�e�~ �֜юX�&��:Lpb�,�LrXI	����N�@�� 1H@W?�9G�~��d�M�$0�V�L����'+�f�f`���=+]Ԍ	�L(QUQ`}���ɓ3$�3~d�I0�̓�L��߫�wt�(���X��2]t?�,B�y��<8�n�N�<��ǲݹ���ml<�8^���9Gn��&�T�u�zl�0�p���,�NW ����Iڱ;I�-7vfN���3���{���wR�>�3n�AO�%"R%4� ��?��?��6�`ڷJ�&pH��� 쓕�;�٘�px�/��I�����)���T�fm��:P�$�2M(1v
��iF ��s~����__�(����M�ll�'\;�3 �\8{�e�l�p�1��2��@�On"����pg��3�]�Z�ݞ(���*X˄V�I�.�]�lM*o0	5Àg��^&�W ����=%8Zh�� ٚ3Vkw*��7��ԩ�����v�*�n���:P�Y�n��&(�����7siP}��g�fI���~8w_�^ wnD�I;MPS�m�~a�$&&C0�{w����‿y�x���3�+Wq��X�I7I�����3�r^&�p��3 ���i�}�&fg�H�	u�t䳧I�:�������a�'b�:!��bC���i���;�T�;ƣ�����C�Hxq;4�ܙT�16�!��$��Lqں0��y�"��m�Yt�C��t��.�Vh!=<::!�	�&��8u��HMä��62�3�f�#~�t���i9��/RIҊ�jKWB��-Kŗڑ�1�� pl^�l  @ �����&Rm�rR�u%�m�ꉷ9Ԭ�M�;	�R�Aj�����ZnGX�pZ�ak4<d��ӷ
W�� (�b{m�؝)�m�n��� 6�      	z�6H8 I����-�[@ ���� �( ��
P���� H�@m���� �t lm@N� 	1!��-MD�zt�lkf���h����l,�釃��1;��:{p�%�lՍ1{tMo�T+m��#g��UcbOn5���!c��y�G��Z��'"q����z�Y�3m�e+l�qڡ���[������B=���f�M2"�����'Z�U2��;��gn��<=s��A6�����.�ۦ���B�U����4Bp/��yJzY�pq%m\N��l`��i.��X���Mkl�����p�0iݻS�VD]�']-��*�{=�8 �擓�	ɮ���u��u���W\�,cP%���ٲ]Rݶ�iđ�����j�u�ez�ֶ�ɥչ�T�J�QҘV� 5�GU�R&(��8�1�i��y�����N26�
�Ie{(�P�Q�@ul�9�B���A�0N�N����2�2aya��j�c6�/N��K��m�N��'���.T���E�ᶰ��$���� )�˫7bM�t���c��H�s�<>���emd���g�9e�e�uζN]����˼Ηs�:�Nʆ��䈱�Uns�.�j6{\����::��^�f\�R��k'��c�c�P�m� �U��v�  ��g��ϋm��ݵ��\��ZY��ӝm#YE�;R�h���,� G`⪅�mR�+�+s�7<g�Z曞�<�8�.5Z��5��Zkrs����Z�:z��jXM96��U\�)[S����n�t4�K�+WJ�5!��{]I���}w 	� J@>��x�v��b8(`'b���Ý]Yۅ{�zØ�Y*:�:�:��v�k�͚�������.�T� �]u993Œy�kAD������ɲ�Ƹ9�&�"v_(�;��۞3\�5�3<�s0�]m�2N0F���Ҙ��g[]<�[dz��YSp&n�sɭ�q�X��gx�&nT6y���.��Yl�/i�%h�]����9�8x�Cٮ@���i��b�6;Y�w-��7����Zٙ�l�@�U|�Y��Փ�WT�Cc�m��x�Zx��ݎ89u�t�N��g���b������V�n"$�7vs^��ͥ@}��mr�@��;�x�=��u5CB��IN;�S������m��:P��u��d̓��}*����hl�'\���`k�_��	���{�������P��Wj�J������3�r^&�W �wf`����g�j�Z�E�p����I���;�٘���=�ڽ�5��HLm�ưj�l������5�x�E۞ˋT�rEd��N.%�U$��6�ȅ-ի�������T�fm��:~fI������{ ����Qİ)P�*���Ϻ� ���2��3|@�J�}���=�;�`n��M�0��Çۿ|�ݤ��I&�4� �����3�r^$p��f���˲�Xۻv�]�n�w�K�$�����$R_ ��S���*Mue�9��$� �Bf=�޿���/�N��}}}�V�� V$C��ŷ��6�{g\��*ؒ"�0N�u��7^1�W8����i������}�0�c��9/ �G<zJT4+lM*�`��Ϩ��U��k���&��8{홀zG�m���έU������u��Δ[/��ߘvN�$`�6,Č�������uU��M����vP�BaB����{d��:��=�� ���$�c�@�36�~� �?�������O�Se�p��f {v>���xv8p��"L-U��9T��G�O�t����d��Ϸb�h.���w65��e
Vm����o������zw^��6t��f!8{ݽv�~���V�4;N�6����U�����@{ݽv�͚��N��T�(�$��U=��l�@}��ݜɓ���4�_�^��Jn��h6p+�d3$B{;��3w����N��Ra:T6)�� �ϵ��*��~4[X��4�y�ݏ�UW������?���L��УT�l�iYGm�w4k\�rq�UK�\��\��gs� ^���m���m�j�?&��Z���|�^�`��@}��m2��&C0����@o,N�wʊ�R���>,�8{�3 =� �W�X	 Qt��V�YM���>�۷`�٠f\�0$$�g��;�����p��Gv�v�۴��;O0ٛ4�u��Δ�$�ۛ�X|ۿ�˥n�C���i���%����;�߹�}�L�`�V��[V��A5٘e!ee�i51����rS1�Ѥ�:
�$� �Ѭ�Z3X@�퀡QI��ou���m\m(�r�g��Z��(�-�:��uUUIʙJ�v�2s�%���nք��Bn�<�N�B��N�9��_eq��uٲ�Fm��%r[�N$��gd�v'����vȗ^��	���	���rv0d'l�����켧U�=aͧ��Xݛ��bBt�Y#�xݰv#]�=�qӸ
N��{j�@�q�r�v�����u6����^��ww����r|��J9��^9��P�7p)lv9�Tg�{u�(絉�� ,b{K���g&"�����U>����۰nl���װ2�r�MݺMX��Bl��� ��4�zw^��l�_ĒN�a��*��0�.������>�Ӻ�~a�&Nn��8��}��p��g�CZ���|���z8p��f {�>��N�n��L(Q3sO`{�:P�07�{~�� ����;�9/ ښ�lum��q�TV՘헕=s�=ny�ӱ[����vM��"�&����h�;R����w���`�#��{�Àg��;���,�ww"�s� ���fR]T��$$*�)I&=�f�,\�A����3d�`iC
ha���������g���ܞ(����~��T�=���ƭ�r�.!�$�=��=�(����gu�gt����:b�!����9x�8{�3 =� �|���Jn�lt��̔�{v��2L���@{�=�`}��6�_�я��:�V֥E�<��-��8�>(�r�ʶ#k�[v�'mӧ���s��[j��X�� ���{�%���p��f�,����J�*�����u�{'Jｻv��f��I�ym]��]l�IRo/ ����;�I�Z:D�}A�d��;!,HI��$�JfWf_�4�����4a��( S.�%�L��gw��>���x}�=�Qݤ����䇉� �ٳ@~L��7�����ޥ@_��v�L݆�. �DLD�L,cv�O"g�a�:i�$�I�3��s �ar� �vTڻv���o ���^��iP�n�$�/�f��f���b�RC҉xN;�S�{6�jK�����`��ɀs��x�_��F��dR'ai� �{��l|�ײ��g+�vzJT5Wv��`�i���c�����]���9_��N�Q�S���&C�;��]���?����g�B�	��7�;�ٕ�{vr�{�f wv>�]�����ڷ5& aȵqs���W�^q�g�8����r^��=����Qۋi疓i������3ޓ0����ve`�`Ql.�ӠE6[u�2n���I@ɜ=��@o�zՁ�ͥ@{��;�����%i�i� wd|{�2�n�W ɻ3 ��r���Nݎ��(��3ٶ�fm*�snÒN�!�HoF�E��`:lSJHzQ/	��iXݜ�&����.'���wu����;~5��܏�+�Q�q����s��}[�*��r��X��0�y�j�Y�ƒ֎�ۓ;kӲiіu�7b�"%˵��^^.z�<�j����6Ȕ�����\����(�r����k���dږ�h0c(g��GcO68�q��n{t�e��h���:�%�x�'^�N��֣?޾?x>{-����5�.b���fx�M\���s0.�������ѷ|/�.�m[ �pm�y���ݣ�q��Ka�v�F��J�=�K��>x{Av��g���/��~�vϛ�@n�m�ٛJ��=�lw�m��Q\�s�ﾙ��!"����֬��T����BI;��<L<LK<
�N�3@wv��ۛJ������w�껽�E[�RT�O+ ��Ҡ7sv�n��C	����`ߏ����,��N��&`~�p	6L��g+�l�W��)Ziz���ݗn7\⬚���;x��\���EVQhn�$��"ݖ�`~�p	6L��g+�I�fے�݁j�W{͖�f��U����G\��$	�7�$��!!1fuu*�������W�fL����`:,SJHzQ/	�&iX����$�3 ��I�e`���Mݴ��]�i� �d�o�.&����	Fv���7�;�%�%�N��� ��I���=6r��&`�W$������m���:���n\�\�8M�b���z�r:�1�P60ĳ���O11`woW�6���3 ��w�껽��j�%I%�0nm*�$���wou����mi�L����0��̎8�G�Tv�]���آ�|�3<y/���M;9n#�:Chv�i�L�g:�qx��F�y�+xh%�XF��"�<m�v�q�i"xC�٣��5F'�I󤌷�]z��TFÝ$zt��秽�bx�܍�+�X֙�{���xt�'!���p淧����\X�X�\a���50�&��V�vk59��#*<t���Y���Ɔ��K1���4Y�Q��f$�����:�0���]bw�ْ�8rrr���k�3��M�̫	��f��hӮ��v��O}��tv1fa�#Hi(�{S��8CLh��f��asi����P0�b��tl��3��d�D�3��ehrf���O�g���ًKg]��6t�p��S�Oa�w���j��h֓��n��`�	��]�C� zP�BC�|ڃĔP< |Q�}G�;M! !�8��N z�8��!УЏ���"iUG��D] P>�]�{uW~}��U����6ն��%n�O0�H��9���ͥA�	�0��{��<�����4�ۡҴ� �g!�M�&ɖ��b��ɒf��Ӿ�xr&��3ݡ���F�<��l�5�h�C�j���7[�j��Zm})򘯔���O�:�?��l�_�\w��`������M:S)���Uy�ۿ�Ɇ0Ü���g>0	6r��l�w(vӷE���y�K� ������3}�0H�]�O��.�:��5�3}��&�p�f݄�$˚	0�:{z(��w�q!2�Dʙ��,ܝ(ə7ۛ�t������C �d���SV�X�M���1jݎ�8��v���]��^G���M�8�M� p-7Q�`�o��\ظo���$���+��I�1��f�}͊�L�'�a�9�ޯ�����8o�f��r���ƓV�t�k�f�fV&�p�l�\ظ݈#)��Iګ�+ �\8��۰5�6(8BHBL�vo|�~}GΆ[M:M��ݶp{휬\ظ_y��U����.���T��N�I�E���SF��#�630��֮}�{�jU�3Z��-�R\d7�73�k�Y8:�����0Pl�9}u��gw*�-�u%q��]k�M�$��Zf�#X���:U�B-�=�E.U����]�\��8{�sô��TW2U��Ѯ�v�v�+��2�$c�����jl������G|=[ݱ�so6�-mgq�౨��g0�mҝ[�u�\gF��m��;�cn�Q�${T�$�O3!.��X����D;{u��όke���gR���C0���nB�]j�?[o˟E�2{fV&�p�f��I���ӧVզ�Ol��$���˰5�6+��&I;�Ů���BeD�M<�����l�\ظOI���J�J���T�g �{f`���2zr���7ۤwv�M�K��Q37`k�lPę'��7�o�����p��f6]���!��Cc�u+��t���C��nF;X��q׷=/�͕��U�V��Li[j�J�\'�!�M�Ҁ�{6�&M�>wE���b�T[�rն\�8۳�"K�Q���02L�(���^���ߵ�/}���t�&C0̑���~�H��e��%۽��n��$̝���� �G��'�e+�C����I��`|�'���>������Ҁ�{6�n����%�%J��ﶴ�_�0�$�v��73z�n��X�4u*��$&6�cX5u�ɷ��A�Nm��=���7-�7C\g[�׷@Q��˫���[o��Ҁ��۰5���5�}�=�`�9�P���H�12P��w̓;��������N�ɒ�$�BMwo��ZV۷uv'n��������$X>ɖ� ��d���7̙�Z���>�(}��`|����ē�D������&�{�,ݞ({3nÙ?FwE���b�TC҉xN���&� ��f`�"��$Xm��{����������R��H��d��۫�3���E6�.[����t ce�{��{�wo~O��c���N�t]ݶ`}��`���7v?33/�;vx�;C9C�!�����%�EϿ~��;�}��>��p�vf�J��O��t�մ�\���N�~fv��޻�;���j]ܖQl���o� ���ݗ`k�v(6��y��O��� �i�M*-ۿ���g �f`�"��,n�px�0H-��hI+n�p-�>�ض���&�r�4T�#�aeF��܂��9K�)���]�m�U�'n�΁���.�["�=5Àw}�0ܗ.�Lj���;���,ۮ�홀wT��;�a�O����0�̾�߱`�l������"�6�R��ݴӦ�w�T���۰>��z�=����ep�7�w��ct464� �נ/#۱`}����sn��ff�c5=��l�0;)f�=��^���i%�x j��![.�T睪�{"g�M�N����.��������7�2��Dݲ�ù˵�x�N1�X(#�7+���G��=]�;N��+��ѻG.wkq��p�4�	�J������S���m�江�N����̯n1�Xx|m��e��a[kmcpJ<c^;nշm�Y�׷������jms�{���Ol�6�q/�m�w4k\�rq�,U�]�k��ܝ���O9�t�
�≦�QQ�D�r>��_ߟ,����;�f~���_ �]ܖ�j����,����;�f`ղ��zE�����ҡ�j�Lm� �͙�wV���� �7��;��6�)]&��� �=��,��_�ٳ0�IeZcWj��VӾ�^ذ��|6l� ��|w}����iU���;��K�l��<�\v9cU��X+���s��q���ξl��5a��,��_ �͙�ݏ�{W�X��(M��v�7E�Ӿݛ36��vH�
0'�ڃ���V��϶��܍݋�נ=��b��m����؛� ��|ڽ"��&w�����޻ٲ�:w����C�m����[/�vM��~�;� �]���5V��k��;�e��٘����zE�J�1շv�8�*+՝�^T�q��ö�;��-��v6s�2;q7!5�[��p�<���� ��|ڽ"�퇯e�7��;��6�t�V�� �0;��Հv-��>�ͻ�N���!�D��LL��L����`}���`�	�C!�����$�%��5>]�݀{3f����6�*K�'j�8�ŀwV��ٳ0���9�3��wE�����T;̼(�C�17�;�f`wc����[/�f�����]]��I�D��|�=y'��
yd6�-�h�ɻVGq�����B�U�]��&� ;� ��H���|�6f��/�Mܢ�qEm�&�}����ݛ3 ;� �]ܖ�j�S�1s5��@}��vrd����M�o�, ���N�]��۾ݛ.�>�٠=��ذt�!�������4hBV	@��ي���s���}V��EZUm+I� wv>�^ذ�pٳ0	�Dpt4VW�ac�:y&{��!p�a���2(dv�l���v�nY5�ͷ��� �;�f`vG�3�a�q�u|��U�8�j�|�6f wd|ڽ�`{�i���Rn�-�|6l� ����zE�{uÀOW��R�[�'E�lM� wd|ڽ"�=�:Prd�������ҹBw�a�L��w�=��,=�e��٘uI|���8C|>i�.��&�(�&E�SR&s[(4l�d��-Y�5�|Èo{f�xY����#��c���;�4�t��,m��'P�a&��ٙ� �Ɋc��j�f�`%�f�\]l&�lB�q�
���M	����	4�{����c�͒Ĝ�ۉ�������b�    � ��ձ˦��%�Z�j���S��b�L�B�\�s�@����3�zqq��]���vyNN�/@�O=ZK<X2C��ӆm�t�`-��l8 �`      %����8 I���lm�  ���E  m�@����� ��A�mpn��Y T� ~�|�t��� ��������mUW���尝�G7W�z��g�l��2\�ljݏ<�pm7e��+�g�fs�����<a��O��]9 Dv�ӌ]�f�n��V�1(j��V^�VI��33��#җf�9{um��v�a�ӌY��뇳��PtF+m�6���䰬�Y:�3�K���i�t]sȖ��	�N�3�ݶ��r�V�M�Λ`#�-��[��(�GZ֫FK [i6kkgq��z�m����޽����T����1E@��p^ �x�c�blV;R�(�Dn��n�"�pa�n��]`0���gn��8�1DFh"{[�����/!�Z���h=d�L1��;\��0[�6s�����M��1n00�^�Wu��G@�@��x�OXv������En���Al���Z�ݱU��rҲۃ��+�,o�N����e�a��j�v�l��7�v�+{$�gc8��g�9�ܸ��A��\����r��n���J��sj�Eꭀ�mNݠZ�Jg�g2�\�vۖ��\��ݧv� �b�G�
�xW��ʽd���dT}��h��Ԑ�`��P��T�;��Y�Ke5�pk%��/n�n�u��vp�B�7b���ٱ���6܅��=�<���S�lۛ�3�99^��ű�h�1�kC�mҜvʷ�Jq��H��ϖ�.��7Z�:����u������y�����p�Mr���v��IH��z8C�Mn�r#t�N��]]l-ӄ�֜5�U� %3�Es�t��V��F��4Z7�oz��`� ��@�	���O²���6 t,� � v�^��׸���O�hf ��Έ�r�is�����	�����m:�E`���r�2lS����ºp�Z��g"�V���Oz������t���I���>�H9«��k9�gl�u��g�6��[y�fOe��Y�צ�T�N��lk#-2y�"�0d�i�l��;��ù���]�k����^l�+�(�p`w�q�]v�8-�^��d�mY+\����*Ij�UIu*��)��a �Ilm��"���뗹^�y����ף��LꗰwnM�6�T���5V��k��.���|�6f�R_ ��H���P]:@Һe	���ٳ0��%�j� ����7������U��'�uI|ڽ"�=�e��٘n����1��M�l����[/�wf��?wc� ����U��H��|X�'J���������=�<P��ذ�ߓ�Pa 28��0M0~m&n6��㙋'g��h�܀�w�>.������w�,�����6t�3#ٱ�&I�p�� �տ+��Z�HN��շ�v=(d�2=��'J��۾I�vs;�r��,��C�LĔ�gtX̝(�٘v8p����`[��7Mc|X�\8vl��8�zE�݀O򦕳�۾ݛ3 ؤ��^�`��$6��aj�-���N[
�݇��Js�j�;��a7�P8���ʊ�ߨ��r�P�i$��V���I|ڽ"�6)/�wf��;u$�i�.���I;����I|�6f�n�rI�Ͻ�D�t�L@�QU�w=��m�jFS�3�@�Jt�3������b;s)ģZ�5 �$�i%H��&��B,vf��F9
x!�(x׹���lX��R��i�n�-�|���ɳ0�Àn�H��ÀOW��R�[���66��v8p��&̜�����ݻ �͒`Pn������C�s˶��q��q���6k"G�[����u�b���[ǋ%�V���~�۱`{vt�>�wo��̾w��~����Yl�T�5��`�K��0���=�6, � Ӥ&�����vI��p��褾��*����[hI��8��������}�r��ڑ؀`ȑSa8���p#H�:u���0�
T)*BRI(LJZ!Rti�t$:�R:A�a�@������6��
ʴ�]�V��n���ŀz)/�{�L�7d�pl.�eYg	r��ݡ�1��F�<��d�6���"�Ԣwiw$ Zr�NLO���2e�E%�vI�윮�)�`�T�i�7m�j�-�|ݒf�8��ŀz)/�_��=ڕj��	���݁����F�Ŝ̓�tw=����=#�J����H�M���)�`T��=�&`d�p���e"ح��M�X�5I|ݒf68py}�����A�4��,D,��I% ^<�+�l��u��Z���7e��2H<��{4q�%��:� 6Zp[�ܶG��-��Q,���.ԛU΄�G�7V����x�����@�	:���iu�t7�S�k%Zl���ܽd��&���
 ktnq]p�b�um�g����.;>��R\i���:�Y:#+ly�b�ȅ�5[lۊ�YoG^II���%��Y����A#v�iS�녑��Z��&e���:G=����&�o\ ���du]��7Y���M��<�ݗ]Ύ�_���`�i&~6������&��@{�����/�;c����r�<̼A1!7`nl�\�L�;����`}�_ �d��v�d�i���MZL��� &��{$�lp���r��WW��t��>q`��>�ɷ`nl�A�$����`s��(x�/2�a13@}��݁əv�q`fFwF M����1�t�ڻ��bv�]��{ocn���m��Y�9����C�\.Q"��'V��IЛm�68pyzE�d|��f펥*���?4�t�l�^y�>�]`	ĥ�^��҈VW���#��&`T��6z�͔�b���7Mc|X6G�;�&a���Uw���pտ|�d�N��&ꄆ���0	�À{��,�d|{���am�HV������>��yϾ] �}�����l�'��+9P���#3��i�ݳ�v7SnlD�.׷[;n���V*����	��%MZL��� M����3 �8��=��"È�t��>q`� ｳ0	�ÀgV�Y�UW몫>���l��E����f���:P�(fd�Ʉ�|���~�^[Ȱ�G�'k�]�V��M�lcO0���3�v, �#��l������(��+t�l�ջ�2d���`}�޻sgJ��e���xvyٮ|���`7k6��ۈ�5�gD^/)����`���.�'i!�l�V8ӵ K��.�}>���f68p��ŀm� .�!ݦ�N�|;홀n��^ذ�G�7�YR�am�e�Ly�n��^ذ(����3�٘Z�H��6�Kwp���HUO��ދ;��{6�-���3���C���V��=�٭�r�~��W'�����t��7ŀzG��3 ݓ��;��T__��4��l�֬�[sw{i�	��]u@.и��,zK]��E�����tۢ˶��>�0�9\�[�`�ÀNע�R�[���62��vNW?�-ذH��3�&`��*��͊�4Ӯ�-ذH��3�&`�r�Iwd��ݍUڧV�>q`�P��0�9\�[�`r@.�Hwi��؛8{d�3v���3b���Ҡ<�2M�X=��^����6��ݥ�%���t����	%�^ 6��vU�(96A:��ɞ��6ֽ���ut͐��Q������Q�y�<z��x��%���rm���3�rmR����a�`�H��u�K���\Yjۂ(��@BV!J�.� {C1vl���e��<.�k��cl�pg��e3YM�cmYl��r�b^E�PM��l�����U.�%���w|����e�n1�r�E��[�}[�gx�$��Vv������y�4�8��t��-�4�0I�+�w���'+�gvL�;u$�`�]ڦ�n�|�b���;��Ԩ�{���ݥ\̙�;���
抡Bz��Õ3Q`wwR�/ۻv�9\�[�`���`�N�t]ݧ\ߌ��0	$�pynŀI'+�Nץ+�)�lcy�I'+�{�v,I9\=6fʹ�F�[L��ݷidֹ��5��k���v�z����k�<e����EM�!E��K��o�~x��,���ww����"9d�;[3Z�|溫���:��,BL�2JbZfb ��Aٕ�>�M���ذ\�b�N��uE�Q*��nm������ދ�����������bI����I3?wu� �)>X�9\=6f۩ ���-Sm7\�[�`�NW �M��l���$6(�e�$�M�-*�S�I�K�l��>R�.�^�.�2��0Ƹ8�d8�d����R�"��Ï�X�9\��3 �'+�{�dX�D�$�6Ӧ�]�\��3 �'+�{�dX�9\z�)]�H�`���d��a���'���u%ٛc���E�ZB@�x����`fw��F:�B�`��q-W�;6��&C�du����.��V����g�d:��uC�Jkl���\��5���mk�3FI�XRPR��%��yhM��N|kXt����	��J��fŉ.��z�ߺ�5�`6�5xoE"�(�Ǜ3����f�}��N���4Nk�	-� ,3}(i���X&�v�!9�nt�	:��ln�mjgV)�i�on�٢bӡѢe�t3���!�/�ꁺ�N�j�7}�p<�����0��kh���x����)�!�����
���N9�^��K�i���P|��v(h dL8��!��ؽ/�*H����	2�	2��3'���@f{6�n˚�;̈R��TLĪf|��s��}���٘�9\�]�{(VӵV�դ����r�}6f�'+�{����"%M&�M%i6�62��T�8��;g�F+yG�>���n����v�����QhI� ���7d�pw\��zI���,�M$]����d������r�}6f۩ ����M�n���K�=$�p�l�3v����i�*�K��T��v���6���Td��rq�:t�H����Sj���y�y�_����ԓ`�N�tYv�p�l�vNW ��;�`{wiP̖���<��/�%�;3ɜS��G	��w4g�4��F��/	Ѧ�~�]�H�&&�&��$��W �rw^�����̒�go]����r�.�t[�I4�{���NW ���37iW$�ɝ�w:w7��$'�)�"����@}�ͻ3v��w^�˛
-��m�]�'\��3 ݓ��=�$X�����d�&�]�ci��'+�{�H�I9\ޛ3 �J*���}�?���\m\m���	9���e{a�]<s:��μ 5V�v�ZI �2s�	��n׍����k���w.�����&�Dql^8�cύ�g��l��b�	�CՀ^�	�����%n�3c�;���凗Y��Ì���n�m�N0�lv�:N9Gsn�n�Cj1e��P���sF���.��ck�^�j�nX�]u�N�u=<������vs:���#+Ӱ���<��3�a'p��阍�����]$8G��::��6�-Qb��7^E��,�NW �ۛvf�*=�Z�T(U��ª�,n�*��۰37iP�7v/�$�a��_RM�m:m�e�u�7~�f��J�d�����`gwR�=��C�j�U�iM��'+�{�H�I9\ޛ3 ��)R��Wn�Zi� �T�`�r��6f�'+�g������9�.u�������8pwK!v�{��zSvxܦ�k��t���K]��_����ݥ@{ۛvf�.J�3���`k���P仢fRw�"U�nm��!38�d�P��+�$����ʜ��@wG�b���Ҡ3�hl�6�v퍧�윮�"���w�}�+�n�>��RAP�����puI�'+�{�f`�r��2��(P�/#�UTX��T���`n����, �Vܕj����m��'�I��Gv6�����َ�7kr��q�����K�m�m�M�,�N�ߧـn�����p��+�{M��Ԥ:�E�`��`�Àz���;�������=#�JT��)մ��8�l\����p��5$DD֓2J�&ęS&VfO���N�ۯZ�q��n�N�e��NW �wf`�:P~I�|�ފsD�C�Uv��pww��7c� �͋�wwy\~>z��ݡ6Iv�����C�O�ݞx8�s�m�-Gs�{g&��������m�2�O0�Àz���=�������;u$�An�V7i3�z��ϩ$����Ҡ3۽vfΕ̙$����\�(OM/#�SQ`gwR�=�fݜ��{�����1}���d&f%L���U�:���T�sb��.d��!��d��J�7Ԩ�6!�5A*]6M�6NW �͋�o�y\�ݙ�lcG��ӻ�m&�Ӣ�[��<;[;�3�	���ʇV:�v]<%ngd���%qN����u�=sb���W �wf`d�p�u�M&�T��_�&������l��� �ﴫ�T��U�ZN���3 �'+�z���7۸�����dM�	.s��J�������@g�)P�3���׷HCi�Lv��� �n����`nnҠ%$���%�FD �胨+�%�\󹼝��n�漝7�ר �kp%��0�y�*�gj��Λ���ҥu��FYĎ#�����[�
���.z�m5ў.[�rd��]�Hl�%q:-u�]fӷc������޶�X��Wh>Q����u����Μ��*��(��B1�⃁|�JN5�%%vWG�Y�t�=�kd�96�l��Q������K���W$��>�U��$�1�1Lƒ�g�,`��=Mrwl����6��P.���Kz�q�_<�>po�����J��{6���Tnm* ό�WiնӦ�e�\�홀M���6l�p��+�M�J�JC�TZ[V�X�����T~N�����޻3f�)R��M&�m���UUϧ�\l�������p��u�M&�T���V�'+�{}�0H��6l�pz�f���R�An;baQ6��=����0t�8��N6�@�N
�nC=�V���qͿ�ui:��l��8p�9\�ק ��d�[v�v����8q"Y�D;P�*�߹�U߾zpwvfۯl�C�V��m&pM���kӀ{��0H��7}fִES�O�R�14�9�2}ޮ(��ـzG鳕�wmm$�6Ӥ�;��%�6�fe��Ł��J���}�o���~�-)�@H�0���c��v���؞��օ�OD��t瓮���:PnuV�i�bo0lp��9\�ק �wf`c�JT���ZN�i�pM���kӀ{��0lp���R.1LD�!Jx&-X͝(}��f3/&���Vd��$�H+,`c�1A*�uJ�/�R���:`��b�:����B����M��ݙ�{c� ������8�� D���ݴ����8��W ���=�٘�tN0e�Ꜩly����KO�7c�t�k���F^݃�t����T¤Ko�o����*�d�@{�ͻٳ���2��*�Jx$u0�J��l�\�w3۽voO�{�� {G��`�%�r&�r��3 ��鳕�;�zp	��[ƨ%<D<L$L݇2fO�����K�w���g)h��d��>� �I���PĐ�9���B�͖E(���*CzO���ۀz �J�`R�۵M6�鳕�;��W �wf`���7���h;5�����ѻY��{qƴ�5�v���nܻ�4b.$ڎ���h�q[���\:~��m��9\�ݙ�{c� �����_��T�"u3,D��fm�$�w3zx�3��P{2�k3's�8:de�q�$���7��ۛJ��ٔ�}��`v�Ic��.ۦؘ�g��W�O���v�｝v��̙�z��71ͮh��R����14���T�fL�ٽ�U���7W^��U��������TUW?�������>�U?۫�&ZR���TPԀ����`��"*	����ڪ��@f`�����[�'��/���������_���~�����+��_�������?��������������������EEUx*���#������~����?����**���������v}����0�����?�?��U!A!D� �!D�Q)Q"U�D�TI%D�D�DI$�%D�%D�$Q%�	Q)dQ$�RHQ)Q(Q)h
B	`!�"BI@����$%`d$d $	HXIBB	XBA��$$d ��a@�� $IA��d	����%$!a	YP��$	VA%	��dD��YE�!RQ$P� $I���%!Y	V@�a � 	YR@�F%`d �$�&� �P�B@�%HBD�$e	@�� � �& ��@��)�)F@�$!
 �F	a�&@�F	a	�i!�a�$ 	Q� YFF ��e 	XB�dHBedd?�H`�2*���2 B� �,#2 ���
 , 2����2�#��*	 B
�����"� �2(�,#0��B2H2�(����# � @��*��"J2��H�0� ��*�2��!*� � �0*2���@���! �
��$�
	(����� ���� ��#	��@�����!"�� J@�� H0,	� B�� @�0��I(2�	�B���A(�B�!)(��!���0�$�CJ$�, @J% ��)�)"�$ J�����
D�HB�),"H@�,
D��"��$J%  ���������"���������]������]������罚���W�s�����O�EU}�G�?���}�ǰ����QQU_�?����䊊�����Ҁ������3�۳��o���0٧�1���4pت*��������TUW����|zu�������#�F
�������EU�����?���Q�������������<��#���TUW��v{��l�_�w��G���?䊊�����0�6�����s�/u���������G������)��T��	c��8(���0�7�   � �t(  �)�)�         
 O��� @B     �T�
I	RR�*��
J�"�%
�(��*�B�(P
�
D�    `@%    -M}���W�8��NMz��,���|�}�vx�>��t�Y\��Wq��������� 8�lf 3>�
8'&��:�� �GՏ��R��к5=7,�c�  >>=   d� h<,��9 � ��= �  K� �  �  �  �$� @
 D � 
  5�� 0   tX��ӤA��g@�B��@@ '` i Q�  è@@ �   h� D  G�xޕv�y׻�<� �����������]�ۏg��w�goq����������  6�&W[�wOY�> 7�J��;n;;�O;;f�s�;k�@��ϓ���ƽ㜼Y�'u�������

   d (��s{%Ɏ�rҪ�z�x Q��m�����v�}c�}�OJg�L�}޷�7�yۯ  �x��8��m�=�Y��q��{j�a^�2��AI���g�����r��y<�٭��D^� 
 @F�h��Yj�G׋����r,�rSw����發`���40 ���ˋ����x  7<c^��-/N���ʯs>^�<����ە��&��>@I�<���׌��Y\/x�t��    i�
�)   E?�56U*j���h"x�T��   ت�=)5H  )���z���   ���jJ�� 2��/��M�Q����I�Q��2s'�2I�&e~��$WQT��AU��AU�DV ���=�j��M~ Nd��#MK�g��Z!�	�a$X@��.�u���#]���I�L'��K��s|&��%<|8Y]ר�����Z���IK�	cR�k0��
s�f�Ys^��7i
1�:C��A�c<�R&��b2��w�ѣ��w�֡s�r�c�?p�s'=�0�WP��_<ߛu�S�J�0�*��y�'<�H���k��%+	���SI@���2n��&>y�n@�ћ�'0� A�4bl�ąd�f�������i�]0%љ��$X�9�h��ښ��a�=�Iu�j1�HF0�^h��c��4i�d��� �5���1�6B��JH�$����
]�n��*k�c� h!��3^j��$�� ��JF@���y��rV潛ד�<�������$�M$
������yύa�/�&�M!3��יϊx@��y�ci�y��2Y�4y���3k�3a J���+f��C���8�$)`l!�1����|:}~7Y�_���OO�O��>�Sݼٳy��W�B1��0�
���f�D��t�wL���=����P���2�dd�}2�U�<%4�����f��n�x��	OK�6߈��OE �w��Ca	u��{�4|{,5mcXIr]j��S��i���Y/o���[������wG�{�ь�c0p��sf����ꐇ��h��ϰ��9�>.���|1������C��g�Z����kFУA��F�(�0�D��r��}.]��F>i�; i8;�P7�Z4MH�0�/�����h�IlaR2nπ�{M��q��$t����:��$,��|����h᧜�sA��2�����2��z��M{��BSG�����+�����^���i��.����Mq��<8$��rp��C�Ѿ��(�@"�RT�VL�c�%d���I.d�	�|��CR$�
K=K���`�@��!S^��Q4�۽k�krg�ӣ�
0��5�n��ŨD�-�{oՖ��V�Qs6U:/W�J���h�ׁ"�BB�eSKb�	�_9��Y1��׎��S��P����>H| �gɯ��c���|k�ͅ�1�q�_<���ı�m"�f�"nJ���%w\��<��-�z=��>�s�4y�p�k�h� a'�mM�fy>O%p�Z�~�48{s����H5���F,��Z{ƺ
S�F��fٿy�!�y�9%-�6į�3a��H��6x���mۨ�!�م�i���/y��>�$T�@B� �AFB�*D����XB448�������_��y*�a ��)
�� iHN�M ��*�`������$��k�
���$bI"���!Jd�����u��P�HNO��IF$B$`H%�I�W�F��Gdd�"0$�
��l�Z,�槏�.��!)�Ҽɞ�d`����xfy���k��Oi��4P�q�zݟhɟ!l4�<���I'#aP�!����{�%�����%߄)r�Ա��&��n�t@�$
|��h7���}(ҟ�Ç�	tns~��X��pI%�"��s�8|����7�w�|��rz���>�i BH�)$$�	V%�<��#Zc�l̯����szI!�#`d���<�ɲy&�ֳ�1�I�)�2:}�y�P6��O=O�m-�5�Y[,kM�C FB��YI3a�sQ��FO9���6r3A���>B$sQ��C�!t��feI~�`��lkO�f�U��c�N��Y��7$!1�'�4ϡ�Ò�=Aׄ��0k(�d�p!>d#CC�7hj�q]ɞ�z�/��+�����������*ӉM�E//* N@2D<�y�
0!g��>004�}�OX1��$	&h�d��n;R�q�4�j�I�ɣ1���Cp)u������y���h�I�q6Sa�y&]�(O���C��p�4B�u����.�m�|y����}u��l�0�m})�b�0>%�!�b�Bi�&�Y�k4l�H�aM҄$(�ָBh�G�R��8CD5� ��]@�H8(r
RG�C�P��o�62C�p3%3z�o�81j�u�Fi1g�FxW�|�d���)]
��z�j�㬼�N�]�WP�0��i͟28�Ȑ���k��/�s�$��L3f��taG9�}�P�O��g�4A�,R�$da�
0����� �B�Y4��a$l��d/������F���M�����.���F�UեR2�f�ͬ������^]_�ⲗ���.Fh��Nl ���,B�CBE�c �a!� yn��y���B�$5�@=S��eY4ӏ�1|$]�����i�m���瞞茜�g�)[<��C��g�4k�%%!ș���!@�˲I]����	(I0!(@)R]�ލ�̖f���8��?���7�{�<�p�daaH�I�6&����n���a{(R�C��Ho��k�$����_��u��+iXA��ٿ8o��}�P���a�(ā!����kS&���Cǎy�a�7sZ���6?yO<�6'�&q%b�~���J�)M)����}�<&��u��ńD�M�q��o�=4Kxx�I�F�CϹ=�}����)Zy���.�#�>ѧ����s|7we��qg�ӞC,�xj��!Y��!�^df1��SST��ތ�� Ga0��,=9�}�>��}�9�(h�l��8y���=D]z����*x�	�� h�.�>��$M�B��<��K>0M, H��!>7Nn^��ۺl�0!`�3*j�I���,tsq#! 2��ܬf���!�>!�".�p���B|m$c���kO8G�y%��K&�j։�ּ7/3F�͛��)�h�B�.y�hL�L� Y�F�&�Hc)�v;�f�(��p�u�#> 7��H�`}��M���� 	2��lZ�0��S���G���R!
k+ϓ,���{��>�<����o���̘ٙh�= n�f���g�'2O6�HS������bPщ1�"Hjّ����)	m��	�<,�>`D�{�G����=8B�����M������$$�s��5�6�hu�͡��i���S�OU`�Q$+�8���;��a�ܻ�'�5���T�H�3R���q͖��ƒd�����4Fל�=��X�O��S&o���')��0��O	���5��8z�4�k�x�	�>k ��jy���b��!�h�v��=��������''�5޼=��fFVf�	�p�����0��k�{��y�]@�&�2bA����>�7)��erBA6F��A���g��xXB��n�z*Oq����!�� �`���t�xs�|���e��'ٖ�l��WR댻������_�O0��#���.�}�@�����J�̭a�7�oy��+�=�l����n}粇��Ϝ_6C��M�)
0�h�7�ᷗW���ɩ������u4#$�Q�"�|�!�I2����l`�$8x��g�#�Gq�ӄޣ�l�j]00��F���4@��֌�0$�B@�IM9�pٚ�-3�C/.�l7\�GF���f�Vp(Q ˍ�w� Bٖd�y�Ԏ�Dӄ�{x\f�&f�[$�ȇg5xO�a���~��HBϧ�֒O�Ág��B1`F0�L׻��5X'õ��A�CA�JB��l6G���xrM|�I;	#b��S�xK#L	�L8i��I$���6�SSYtfNi��Oy�7�����!w���5�b0B�8�$�_	�&� ���n�^C���y��-�B�IrG ����7K�r}-<�<��K����0d��dY���y�>%/�+�$]H0"��~�5HY��]M:yYM���Ԏ���pɣ�j�>��a}"<d�a	��j�d��$�<�>��3m��9"�0:��ā @'@�P�A��)�!�{���j�dbH?��z0�0�w�Y���i��@�܁
�%�9&�٭:�!c�l�6T�9��awv2p�tS��*���C�����$xkWdw����c3ae�h��e Ͳ�25��	!+�˛�M�O�
�Ì���&���$������ {u�_0�����D���sZ�	'���P���槆��N�j����t��h��(�׵9��JiN~��@�ļ��qU~��@�HHV���W��=0�����T����s�;�ϸ��zc�ݿ����4��O4xh��s$XK�k[��o<>���n�O�~=K`i���MIA)��	����d���<�	2�{�c ��	CZ2$�������<����y	�5��VI8����M��kn�r�+;ʷ]J��6i�   l    m             ���m& m��v[Q!�    ��`�    |#�      -�   � �>         -��              |  6���g$HH䲲���t�s�P61X�Z���N��I�ڕk�;[n�"^Ft-T��2�mU�E ��m�m3�e�[j�j�k�F�tNʲ�[[VѝP�.�n�J�
�T����Σ�V	VWf�V݇m�j���G�\��J��ce%���<�����C�#��Ζ�Úq-U�ƺ悧r�
 ڔ� �@=R��3Pq���*�U���nݧq�������Y:I&X�����%�Z���if)0c��Mtٮ�������I��n�׉��gHt��� ۴�Z�Wh.����U�YM�y��b6�8'+�įK9���`ݎ����ʺ��<�C�&�"1E��fU��ܲ&٧Ժz�[ـ䳯8p�V��֧Nt�Ua����X�e��`� Xa'6�]����� ��ć/C7�z�i
YWB�V�ZM��j�+�֬��SÚ��W�A��unz�	�[8�v����n8�	�N�u�N���m�8�:f�ɔ��)���R]yn�m�                    8     �n   ��a� �m�     p    �` ��    8    �  >��`[@     �[��M� �          ��    �              �    h     6��  �  	$�ŵ�� ��           H       �               �|�         [@                         �               l   ��8� :�v��Mƭ�[����  �Ά.��2q���Hm��.�v��jr�R�ÐH�
�@UUS����⺍=�yX +��mʽ�V�c U�P!-��:��U��<a��mPe@"��K�8�b�M�Q%��Ie	m�(�iW�U*�֨6؝�ek8,�9�v��� �s��fv
��M>xɻS��bS��P��'YA�ڎa�Z Zm�nm��T�/3�Y�[d��޿^���7]T�-X�]���[q��v_*��J����oiQ�«�/cZ蠝B���]j�!�ѷl�v�vh�V�ge��wE���V݇qnac���gJNR�͕!;m7J�����eX���e9��U�JZ��������ɜI����Z^&^&I�қ��N��ʵ�y�wk��5���z�s�ښ�`-��bX)�N�
����  � 4i}s[�H��86� k8Efyn�V��D� �i�pFqӷ�[�Ėy�l�5t���\�6	J���`+�)vVruѺ��D�j�Z�t��]�$���Kڝ5[P�A�m1�vm��g8���b�6s�Z�duR�Un�R ͫm��-R݈�Bj�I�/l�R�UR��U �ֲ��+�������z�/Zp�-� �fm�l	���_*�A�8�݆�@��8���4۷HMZ�Y��W�{@�r�т*�e�0�e ����s�-,�񢁴��}����m 5�1'BC�b0���b�NB��B��vI�E�Ѱ�֊k�F�WvU���F�R�;U�TJWWR� A[R��,�&���m�&���m�*F��m�v�5�����UT�*����6ܢ�n�~/���m�+j��`6��ڷ[��z�+�G6��Z�*�	8��fy���j��hH�ԳI�l�l-�!�$��m&6��vӢ�HR�d�����^d0+��j"ؗj�YIv����n�4�h�   q �I�հ�h�&[���-��ۆ��jA[^
���UѠC50��[�~|H�\�۱��٪�j��s2�G�Z�bU��9(����@@���om�Wh��Iu�λ`��n���,g�3��0'C"9W�� �����h5��NQm���ː�����GUF�Y�T�X�*�g<�Qu�uT�I-j;#�*������;uv� 8m[��e�M�R�tee�p����l�ǎ:F�A�M��!nm�� p�gl�n��n� ��K�qUH
���0�ʵ*pl�U�J�+��J���m;Z�rEO:*#�j���C��!;r�R˲�'=��ڤZغ����,���s�i2,�mUAP<�(�mF�Y�m���Bv�d�f[��
��  )�T<m��m��fz�x���{�7nP%GӸ����*UU ��G-P�(U).�KhmtR���*������N�j�]�RX[dI�kr�@k�-�n�d��m�`)v�.N����@*��UT������e��Н�P�PVZ��6۱)2��[R����+j�uM�R��R�D
�V�C��]� ��m�#!��1  [ׁ�l@�[p�I$� M��d��\Zņ l��m�8��FZs�AZl�m�M=��8�Q�g�Ъ�T����l�ƒ�]6�"��U��5+�?%��2� *�0@�3۲���v1YyR�խԪ���v�M��=C�W���;� ��e9�H�}�뭩�X-��y�9ҡ�U�V�b�&ڮ����T۳��h�E۶�i����h/Z8��؜���mwM�_�]���R�&f@�l[4��\#<��W[Up��m�i�k��P ��Al���[y/V�%����)�Z�ʵA��[�`����4�!̼ԝ�jC�m�S�<[��ekj��{;s=R����Y����Ygmp�ƃlt�o��u�$��ݩCR��@�V�ųU+������p���WGI)��Iֶ�Y'We�Z�Ԓvt��YPT���1��ژ�`��H�T*� �UHͣ��̩�[m+U<�wm"�ԭڒ&ub��;m�r�vA�Bkd�f�.���h�D��l�5����@�[1p7f;��\�K[U����ʅ���V�mT�.2�[2��sC�md.����N˶��UR�!�n��u����Ke"{K�*�T.[��ʴҬJ����ZlA��D��	C<�+(\h��"���Wf]���%�WFD�n`:�����t/����rV��mui�q��������I�A��ҧ+�W�Pf�K��K�pI9|es�6Wi(p_>Q�/g� ���,v�T@��m��@3�Qp<v� h�W������8�f�J�ÕWT����UF*��n�E�T������;U)��b������&v�U��ŵɣ�*�*�m���S:6�)� �m�n,�Wq��psv��	�I�u�q��+9�{JR�GJ�zD'\�R��J�R��N�ɶ�I��oVC�%n�.�s�59c��v�Y�C�v���k�X��I�N��j�m6��S��rʵ�JKʺc9�$r��l� ��6�x �yk��>]P�.�f�]��l �pk�������؋���� 6�d'���y�V���,� ��������Cm�0����U��h
��n�rD��n�Hq!��  ]4�+�ݺv�p[@k��E���eKAmckP N��e�N�ҫS�2�R��(ʴ $%�]�`X`��ݰ	  �M m�'HH�����9�;Z��P֩VZ֨���,U˽���Z�%UZG���\�`���惩4-�:����خ�ݻeV��iɓ���
Iba��sO�.����.�f]9h
�S@e�L0&�6<b��$�U������U@���^p�  �ԅUKBXP�'*�%N�6��`4P���>b�[fު5�9���7lհ�sv�h���Z���+5����pj����YZ�Om�=e�T�,{��7|>�*���ں^Z��v��j�-r��R7]-[l�=U膞�.݃���$�`J,aUV�C`.�"[��@�P	�t�ͲMVFkV� [p6�@h���ڶ���Umo� 
T m&L�)�����)V�3�-a4[nհf�H��<��p�!=T��j�:js��&���� v6!��A�.Z �i��y��r�ͳi�YZ�4����i��5�d��8���7M�m&'8�`H��5�'��7!�%�[!��Ƞv��Kl�0 �(�%���j�� t�����.��I���T [d�f�L$-3V�l��n�Es�Z䉨��
���$s*N�⫗���HJ�Z� ���΁��R�v�/C�kXI��b@9gKv��F�4�c�V�v�KD�]<[�u\9�M]�*UJ���v��\�պ�?戂���A �GG��� �Ȅ!�Я�DN)�t�qD?ʅ@��O����P4
����J��c��@�8��x����_ߠ��h��Qb�8 '2IHM"z���pSJ�A�����"$� >Q�D=Sd`� M��)�>����4| H��dR=�!��P� D�"�H��"D�B)`"B1B	 �8' �< Ҡ|/=�Q����6��	�Q0D*!v��F�������A����D�B$���x p$	��Ĉ�O4'��TLB@�S��6/���t� ������*x�T�b�)4&�!�6 �6࠱L8
?v����DC�V\��*��D�i��Wh���B0H`�0Oh!�];a<A("��Р:D*A~��|���W�]��bF#���#�=H�'� D��`P��vUA�i#�}�0A.*��6�|�� :AHA � 
? �$�0$	��9�P�	@�t�&�W�0Q�4� �}S�� ��@܀���G`	�")$U���I3	��kY32ۙ� ��D�6��G���j� p  m���N���\4`�0[��s�<�1�VcvǢx��x9�hv�э��ܜ!M���Z$�S��L�u��˼��/n6�:���xA�[�Jec<�<��מ:����r�%` p   	��ăm����,��6��z�� �	   �t��8$׫m� � �h� -�� �`    6�  �e�B�f/l�n̛��J���d�ʉ׊X��-��{pT⸮�g\�4���r^K��[(X�6�}[vza�bk+�y��d��9��z]��03��V۫������u�5��^w4�ԝ�-��yۙB��6]������-�U�Ck"u�b�2�n��7/gfݲ1��-7ou������흎v�-f�1���'v��k�I� r�U[)0Ln7YΤ��Y-�����}/O!�:��:M�yx�:��w8]�q�l���խ�Q�WKn�UT����[p1q�\���uӬV���H0��Ss���l�D+]�j�,��:�:v<ݦ�6Ht	��G=���h5=)����E�k����u:{1�d�ǵ���9v��Ρԓd�=Y��Ӵ\�X۔��h�as��wl�1�x#x�OD3���t\���bm�;ӳ���f1:�%�r�V)'=����fmp=��=��C���9��c�2իk�Wcn����^;bxun�ۮ��<\�T�7FI�]<�n{i��Ag&��;c03��ۢ�0l�]��s��Τ��bAw#h�o]�:K�j��Ő����m�9���z2ݙ��T�c�ݮz�`�i�k�
�k�z\�=h�;=ln�9w,<���G<�����)��=5v��1�	��ր��OfS�kvNy6��6�Zطgsڸ�7yrގ'a-�c)�,��w\s��R�n:�=�L˙�0֍\��5�K���J���8�B�x
�TL��	�T�*�����>P�Q8�I�/�ɒ�(ʽ6�0��M�9f�Y��n�\�^5�Җ���r�<�gkd
�Vv�뱄�Ʈ6;+��C��D4�ˉ�m�����j'��ql���=cJM�غ�FxSsVB��C�0��t3��z�<�页�����g�3���'x�4�7fL��9)X99�;q�۵���0=u����\�n��[ur(�h��j��rx;@ڌ�9�M֥֦�n���-��Mʝ���D��c''g=�嘌x6`��h��$��E�;�5 ����Pܘ��\�Y�tx�1c�ɠr�V�Q�٠uvנ�� �nT�"d���@�I5 �ɈI5�$��j�/x�H��nM��� �٠r�V�Qm�:åxLM�0��@sP2K@z�&��1��o��م��i���:�u��ӹ͹��ē�kG�.�j��y���Bj��0���6�:d����M@;rb nM@8eI���DӋ@�-�O331g���e}O���˷ rj�Ih:�,����Y"�rh]��{l��铽�n�nn������3ȉS)�/o7q 7&�:d���$��v���kodŀǊ#6��+�hE�h��� �m�����B��p�C��X2m�J�m���zN^v�5�4��u�g�AC1��(����o�~�0y㖀�Px�#{VYw3++sl �37Px����9hE�h�Q�&&Ɉ�@�- �oٹ'=׿]�+�~�W�f��{�7$�j�*���b�'��I4>�<]6~����ڀ��- 7&�9�캨�'�R&�Z��޾ՠ�4z�V��u���FH⍤�j�nݡ�B�Lg1��Ξ�<�����+D��a�u�v'<�nd�6��W~Zm�@���hV�4�]M�&I�5�y���Px�:�ɨ<r��Uo\ŀǊ#1�4z�V���4k32gdf� f�� {����L���H�.�f��_j��f��|1 2�B"���>W}Z�x�J�x�8��rhx�$��9h�2j��wW��ds:;,�=c\ty���qn�u�B�R\�!8�tDk/k�.5��c��j��[�7�}��?Z��q}&"H�y<�@����8�]��}�@;m�:>�eXc�fI����̚��c���P�@v�ܸ����mɠ{�ڴ�٠{��h]�� �SE�C	�bP�^%��2hdəz���ll�Ny�~��|��U EHI	Y;�_[@�*���%�Xw��W̵�����C��;���e1Z&ڢ^����������r�(rn��Gmv��ϝ|���k����ў�d 4k�X�HE6�n-��Si/Ha�rigX�	�l��K�N���ҳ縛�|�����@�l�]�Sr=�����"�4'�.���U�hܦ�u��m�\v,�mM�6�n.V#M�j�K�5Zw������~[|??M�Նu	v�QÍ�̐.{'<pP)/L��;k�t�;Fp۴$W=��#qXf�'�@u��P�r��j �;�8∂S	��8h몽��瘑޻����M�YM���6�x�<��n7�s��hol�yl�;�kz{IZx�6��L$qh�j �I��L�v9h\�W3DIO&<x9&�{�f�޻[�9�ڴ��h��*�Nd�6�R<Uq��o+��˦�+�g��=����=Oi{)���E�19���	Ǡw���q�� ������������H(�{�y���^�D) % "$F+"�b���B��S���l�����<�����uW���h�(a2LI�'�vI�_I��\�o`��w���b1c�@�[^�����9��hm�@;̹\MLQ%0��9�缌�RL�y����٠?=�E��Q�$��Ƈ� -=�aˏF*��On���89t�緮غ���N�[�������5�rbۙ5�ثo�ژ���n��7���9~�s@����;�M�����)���I4{n�����g��x�2��̖&_�NF�������>��&�H���uv�4qڴ��h廚.ʞ�����Fܚ_I��5�"�y2b�.�}��[,����f�a�KF}���:���>ԉ�`)�l猨���up$��ɨ� ɓ?}�z�������M`7��A��@�-��;�]z�z��4�\���(��H1=ݤy2b�9��5 �EH�fQǑ�L���ٙ�����3vh�e*	el$�0�fa	2Ʉ$��Hvjf��s���r�D�ڈ�HǠ�@�-��-����{^����\Y&FG�<#K��;�p;�a�p����Wo0�;�����^I;���qL�I�w��h�S@⽯@/m����Ua���BH���fa8V���[�lP�����T�ʞ��70k$ĉ��� ��h��-���w�������1&��1A�ɒw�ݚ/gJ3	Y�~���@�~_kX�1y$�;� ��\srj�əe��rw�@@�����&�H%�׷=�kO��cS�I=Y�n����Я0�*{Lμ�mv��C�_*MՋv� ^;E�zY��7n�l�ٸd�����w�Cg�cyn���W��/]��Зv5��k8�[��e�t-@qGc�P�7��O�����wcF�U��7C6RǶ�Cs�F�oP�b;uF��@�c&x�׸�m�㋧*,a��ɗB:�&��oZ������ֺ{Rstt���g�KZ�lEl��hb��"#�	��c���@]�#3o�����@y��(/2h�N��`�CkG���{��f$_�����@���{ecmLLq�0�&&(/2h�Njg}�'J�sb�9Ӹ��$#�dx�M��W�oƁ���@⽯@/m���ҫ�Nb!$M�@�����u�~~�}~�h��C8���Ʉ@E�dp�u�b��:���[�p�m��(m��r+׹�.����d��!�q^נ���������u<�8a2LQ��q��߳~�$F$d	��B"��$�D�К��ٹ����8�k�=���������@>��� :㘀#sPW-bnb�0&Lrf�oIM��^��{�=�$�n�jI/{ݢX<�/"=�$��jI%{�=�$�n�jI+zm=�$��k�dN,�C$�C�ck���v�G5
휗-�7<�%����f{!�g*\9�]�i�� }��~ߟ��t5$��6���Iv�5$��N���)���9=�$�n�o��K奔��I_��RI+���fy�����_,k�8�qE$��$��ߏ}I$�l��0�6�	RÛ܄������D|JQ�����G2kD5Nk��2@� ��7j�	�!P�R�	u� D:J!5�<ۉ(�L͑�$kP�D`�	��w��M��< 	4���0\q-��8�8:q5�|9L�'��
�u<��<�¯��; ➯&��xp�3(cD%٦4Ұ8k	���Ț�m	hf���"�_���6�fa沼(�P(���<5��J#�F�D��M��Kf�u4:�DMc�X����d&�q	]��7̼�٠I��>!�ctec$���4sֲ!�q5����z��x1N
�-�Dx1�H����"tD8��t��C�@x�'E�OT��sZ\���Ԓ�����{�x��LH��ԒK�ɩ$��l�Ԓ��$�zm=�$�^D����1GQ�5$�����]�t5$��M����]�RH�-�����q�v��]�p���1����aæ�:��v��������jӔ�9���A�=�$�n�jI+ޛO}I$��'ب֭�����-��G�ԷXL�	�ar�����Ԓ;۹5$���{�Is�t7�3�m����CCk�5��!��RH��rjI%yl�Ԓ�n�jI+Λw�����\�p��t=M��������m�߷�7m��=��s��w�)D�@� XU���A���O��ȜD�~�ᛶ����l�HFI�c��Ԓ�n�jI/|��{�I�ܚ�Iw�{�%޵���Ex����ͫ�qn�8�A7[���nz� �w:��<�����#��csշ�����S�RH廓RI+�g�y�fg8�V���K���/q��$=�$�v�MI$�-��Is�n�J���RK�dO/�L�q��I$�-���\훆�����Ԓ\�a�$�}i4�9�ŐNO}I.��-I%y�i�$�n�RI+�g���o-bNaa0N9.���Nr�z��{�d���{��-��u�K�m���0�� ��T�+��{��~��WKʼ��tQ��:a�κy���2�&�:��5��Q��m������UU>��m����Uٍymu4�҉�ٳ���@F���s̿���>��;v��7`�ź��&z�WS�$��n�+lv�Վ��aᮺ���W&r��"uc�R�j�V���c<�t��y���ƍh�n����:ƃr�(�㳍զ�sMc�9<u9��~�w����_��ұ���sm�$g	;��S�W*o`�kp���h�8�lQ�d�;;=F�^D8{Ē]�톤�W��}I.��-I%y�i�%��X�S�Ȥ���W��}I.��-I%y�i�$�n�RIs�we$#$ȼx''���z������Ԓ\�a�$���RK�ѥV5��C!n%�$�:m=�$�[�5$���{�Iu�[Ԓ\��q/C5&$H{�I�rjI/�x����$�n�ޤ��)��Ԓ��v�#~������k<��Es��g��F�H�lŹ��e:��c��:�۵��Ά�� >�ߧ���[�oRIw��{�I�rjI+��I��O$�cy$�Ԓ�}��|��2=m��RT!A�� � �mS{��ٿ'9m���fn�m�Ͼ�s�x�_'��I���DH&ԍ�I/�M��Ԓ9n�ԒJ���%��[Ԓ\�v��q��O�����w�����o��~�{�Iu>��$��M����Webl����ȞE$5$���{�Iu>��$��M�����I%�Z{�ئ$�Ĝ�ɣ���Mծ��K����=��ۮ7��ŗ΄1=b�����k���?ߣ��:m=�	�rjI%yl�Ԓ��I7�bq�I8ޤ����߼�3h��nMI$���O}I.��ޤ��.+�g�<�5&,�/}I#��MI$�{g����2/�����Sz޵������}y�m�y��$�dNdԗ�fx��ߧ���n�ޤ���j�ԗ�y��~�ܚ�K����k��y&#�9'���[�oRI^B��$r�ɩ$��l�Ԓ��k���d[f�%�hwY��%k�۞x�A���-a���-m���T�uѮѫ
R�+�Z��$�[�5$�����]o��I%�wh�&,H׋������w&��W���RK����$�!k�߼��ڮ��$�bn	H'�9�RI/��{�Iu���$��-~��G-ܚ�K�����nL�ǂr{�Iu���$��-~��G>�fn���DЮL�~����5����%�8�d�N7�$�!k�Ԓ9n�ԒJ��{�Iu���$���nDH⍃)c�u���ϡ��5!�S��]k$�Z��tr2e��:�!��m�fۄ���~ o�߻�RI+���%��[ԒW����IU�U��|"$M�G!5$������g�6�[�7�$��>���Iv��y�g��J��SM|�N�9'���n�ޤ�����W�y�l���5$��ߧ���N�&�"&	�#z�J��}I#��5$������<�d�7�$�ۿ	�4�y#^/#$~��G�jI%{�=�$��kz�J��}I/|�3�3�<���L?M
�,��q������5H�6m�I-"&Nܩ0�T�T�T�qK�j� 5UT����D��0�q���%n�u!/EE��|�~n��v{l�:���]̸3�8˶B�5��a���,˅�0���&�M���m \io-�;C:"�gN{TB��&t�p���x���A�R1�r��9�N���'b�Cq�x%<d��ЎI�浩M\˓.
|�>	9������{\Ύ� �X�X�a�N:�.랴�����2�prv���kg��RI.��=�$��kz�J����I|�������nL�ǂr{�Iu���I+�Z��	��RI+���$��RM�X��fH$�z�J��}I#�Rj_fy�co�w��RJ�~z9q\K�FhU��ޛ��}"��*@u���+�>��}����c������ ?<�?g������T��s�O��f7]���g�:ʇl�8(N�x½���N�� ���:~ ��ۗ�~�sb���2(�e-o�������M�DL"$jG�v�׾y���R�)+
DlUh!�&K��#;�P}Ԩ>^Ejgsۓ��ǃ�����=��4�w4��2Mɢ3c���;����y����9�Nf�ؾ�������-e�C������mIF
A�2/q�@��c���7c������(���u����"緕9��a�59��v��U��0�s���즷t�p3�ե�鄘��"�oa���������}N�!D�xy��f(^e*�M� ���͎�?d�Z�����4SC�m�D�h���9�j��x�7�<�əy&Z�b���m*�a�!�$�Bw����������ؠ=y��?�sF�o=��<A*\�.�2<<D�� ̊��ɛ�ow��ݍ�=qj�-���$���$<ݍ=�c��t�cpݔ�C�≘dx��?�g��}Lo�5�����ۚz�V�λV��e�@�w��0���rȜ��/��4A��@_A��2�w&hg�|��<�)�ȼ�H����h�fE˙%�����@�1�� �N�;�I��$����3zx�.���rP��U��HV��@�.�e���=���;�N4H'��y&b����@srM�[��3c��k-z���FL$�Fd��ញ���]l�3��:��gF�@�1F1������w?0��<~��c����8�?�-�v��A��������:a���$�Bw���=q����N�ؠ/6t�;�ڷ�<�"�~d�ژĤMŠw�?~�9 �-�$�I��o�5���}�x�~ߍ�~Z�3��d�ɢ���-�zx	O#ĩP��Uw�@rd��,��|���^Nd��?$!��7�IH��.fYv��,Hԅh�[>O��(k��"$ӭi"n4��q���H��|�K<`���8p4���g��Gd��`�$Є���Cu4:*FT"Đ�8D�)�<7đ��>��24���@�K�}��d�B!�H��2{�"V''5�4�4�)�,I�]J���6�N��Z$8��JaG��7��=�!$͆�7���H�#B��D6Cxat�4�� ��x��uS
A�'�a�OC��l�r��>@��Bs�HZ�B#!�d҅Y ��7�3	%��HFi,	b Hd�$/�l���u�P��
h�IsZ�#��j�齚bNA�tj����4&92��Ma�sn���+��m�փw�5���Eh�ׄ�=;�>��RF�xR@�i������ ]bĆ���k	q�h�D�*a��E7�hm]��^j�-�3Z�'��� 	$Mse�8 @m� 	6�� &�̎��[	�q:^���vǆq��.�����]�=���L0pEgG��������6��Ǘ�����$F�/`}�b�Z�n/EҔR��9��y�Q�Fp��{M�+�;G�l�@�  @������tٶ�Ͷ�   8  ��A�[�  �8�� �A"@6���      �;[�[7l�MF�e|�f �d#A&���]y7�[p��&v^���&�3�k���=��8��<b%��>|�>{�Ol��u�Ò�4k��5u��mn1����5lݶ�N��:t�n'<���j��m�Ps�2'.�Q5���)�uF�h(�s�Ƨ7sw7Ty2c<#��G0�!�0"��'�.&�W6�8@#h�ۃ�+��b�8�9L��(�݀�'e����k5�w=�#�ŵ:��5�X�j݄���z.�u�������
�)��͸�e㵞��[�Jlp��I���E>'��Ƨ]�v��\&���*�EpcX;+�-�(н��Z�6(�^fMjv^�Ӎ�)�u]=c�!�K�d���i�m����V�=,�8��ܛG3�zgN�C\�/�ςa�snX��L��+p���������	�t�礯&��/-�98݋��K�z�cB6��ƺ�)�����;��B�3����';��w[+��*L"��VM���%�\v�Q5����������:�;�6�؝�9�˝��C)�6�;�\=�����;b�˺��f�4O�=�X0��Q ˵�ֱ$6ǧF�Z�$���Kd��$4�{$j
8�GI����a�9F�m���Ρ��l�ŷe����L;�gjmn�z��sl�e�WI:��Λ1#*�l	�(ԍ�4kl�ò��r�7\�'F��=�7jq��㙗�58�e1t�oO�ZH��U�I,�����}��p�c�٬2K)s�Q�4�E�� ���څz
����>��S�x U��w��w������;���ǘ�'iN�T�zv��:�<�t�f���HMD�[J� ���UR�B��p�������܈ܓYD����7/=s�<`֭dcsg	d�Y�c����L�ci�j����ܭ�繛�hm�+e�Z�kN�b��ȼ��5&훞.���ܧ<��#�T���ݺ�*arr��U��u��;����4�>��ǽ���{�~:����������;�݄\�ΠA�u�JL�6��Vɧ�䓿�ws񤧏4Rɑy�t�;�h�v����y�g�-w�Ͼ>I6�҂^8�q��v��<ċ���@�ߖ��;V��Q\KZ�&�Y$Z/n�w�F�N�q���F�����8��]�D�D���A��$�v���܎�?b�Ǡ��2���*�tü?C<I-���/ј�%�|���v�*������F��X	�m�'�xF�7GO8[>��W
]�u�˴�*�J��������>|���aS��qp�����9{w4�Z��ڷ��#�G�~��cx<h��&h�̻ND�,K���NC���Ͳ��:��T�T�&3pG��F d�1VEd�S�O�@�O�X����kiȖ%�bw����Kı=�v�9�
>$e#'t}��;�Jx�/2B�/��D�,K������"X�%����ݧ"X'�#�����;��9ı,O�w��"X�%���[v�칓Z��\�k5��K�?	Q;��~�ӑ,K����v��bX�'��xm9İ?E ��N�߿kiȖ%�b_�ߧ�n���[��Y�]f���bX�'��o�iȖ%�b}���ӑ,Kľw��ӑ,K��]�u��Kı/����ﰗ]����ԥn�Ų-�+�;:���ᣘ�T���h����� ��%�m����u3&�Ȗ%�bw���6��bX�%�w6��bX�'��{���?�D 0�&D�,O߿M�M�"X�%�����%���k5�a��ND�,K�߻�NC���D�K�������bX�'{ٿ�iȖ%�b}���ӑ,K����պ��u�K�-�ͧ"X�%�����iȖ%�b}��}�ND��z�� ,`Q҉�E�E�B�������ӑ,K��_w����bX�'�}�o0��pԷ2Rffӑ,K?�?��(dO�ߧ��iȖ%�bp�r%�bX�׿w[ND�,��h�&(wwK* f[�<�D"93���ɚؒ	"}��bn	"��F=׿w[O�,K�����m9ı,N��u��Kı/{�u��.�����7C�c^{u��'��Uݑ.[��yS�y�M����=Y��%��=�=ߛ�oq������r%�bX��{ͧ"X�%��}����@�bdK�������Kı;���n��˭fCZ��ӑ,K��{�m9��Q5����~�ӑ,K�����ND�,K����iȟ�$X����%���~���Z�,����ND�,K����[ND�,K�w�6��c��5Q?}��v��bX�'���ͧ"X�%��{/Ky�l5�W35�5��K��V,"~����r%�bX�����iȖ%�bw���ND�,Hb$dXAF	�
ՀH�QHJ��'@^�+���L���5��Kı>�Oߙa�9nsXL�ND�,K��ݻND�,K�I������ٴ�%�bX����kiȖ%�bw���ӑ,Kgl)�(�ciɄ!�c&9�lx�I�.��68��ǭs���������i��3Yv��bX�%���m9ı,N��u��Kı;�{�i�`�D�K���w��r%�bX�}���rLո���l����Kı;����ӑ?b1D�K�~��Kı?}��v��bX�%���m9?+QP2q���<�LÂy!䘦_�Oı?w��ND�,K��ݻND�,K���6��bX�'u�Ӻ�r%�bX�k���n��W%�L4L�ND�,�Pc��\���~��ND�,K�~��ͧ"X�%��}��bX��B	������ӑ,K�������f��Y�P�̻ND�,K���6��bX�(~Hȧ��g�m<�bX�'����iȖ%�bw���iȖ%�btO��c��B��Y�~� �n��Uګp�y�u7=!9��|������������z�h�T�P�= �e ��2&�u�;Lh��nj�s:�,��2a�f�+�'���7�x:H^�"� ���P39ř��7jH{F.z��ۭ����Y:��$s�]3���My�gV����9���"xe;c'W���;V��V�+=���l�Ft
Su�X��s��h^�+n�q0�9�c���ܜ�v��ާv�#�q� �ΰ�+s�5shF��F�����q���X�������"X�%�߻�ND�,K��ݻ�W��}��,K�~��ͧ"X�%����_��j��d����d�m9ı,O{���r�`���j%��_w����bX�%�~ͧ"X�%��}��bX�'�'zǙ[�\�Bf��r%�bX�׿w[ND�,K��{�ND��E���D`F(�L���ߧ����bX�'���m9ı,N���[��M�Lut��kiȖ%����A #���~ͧ"X�%��]����"X�%��{�ND�,�@�$SQ?g����"X�%������f��VfKe�ͧ"X�%��}��bX�'��xm9ı,N�߻��"X�%�~��ͧ"X�%����~��L{��nm���8I�=p��=�����GO:&z�3Ԥ!ff����H":�s�SP�P��8'��f)���d�'o�}�Rr%�bX�׽�bX�%���6��H��D�K��ܝ���"X�8��N��%C��$�	�T���ı,K�{��r��>�P0A��2%�w��6��bX�'~��u��Kı=�{�iȟ�P ��j%�����jO�5�Z��]K��ND�,K���fӑ,K���>�c�D2&D�����"X�%�����ND�,K��gm��[�KMfk3iȖ%�bw�w[ND�,K���6��bX�%��m9İ?�c�ș���ٴ�Kı?K�[g52�Z��Ys[ND�,K߻�ND�,K������m=�bX�%�����r%�bX�}�^�iȖ%�by�~�� �ᔱ�f�)�ۍv��ųj�TN�6�u�3��u�/��rDۦk�"X�%�|��ͧ"X�%�}��ͧ"X�%������#�MD�,O����"X�%��㻺����fXj]nfm9ı,K���m9�.�j%���o�m9ı,O�~��iȖ%�b_;�siȖ%�bzw��u�����l����Kı>�;�kiȖ%�b{߻�iȖ<�+�O�P�r&D�����r%�bX��{�6��bX�'~�}��ѫ2尸I�f���K��O��߿�6��bX�%����6��bX�%���6��bXȌ�N��k[ND�,K�v~�e��\�Y0ԗ0�r%�bX�����r%�bX�E �5߿~ͧ�,K��s��kiȖ%�b{߻�iȖ<oq��~����\� �[t��V���:Ϭ�'W��s\!{tm]1��f��kSN�m�E1�r��G%̚�fJ����yı,K߿~ͧ"X�%�����[ND�,K���ND�,K�߻�ND�,K��Ӷ�n��%���5���Kı>�;�ki�#�Q @12&D�;����ӑ,KĿ��fӑ,KĿ{��ӑ?��(����"X��������L�֮eֳZ�r%�bX�����iȖ%�b}���m9ı,K���m9ı,O���Z�r%�bX��N��2������ӑ,K? �`E�D�~��m9ı,K�~ͧ"X�%�����[ND�,����H@jP�H�$"�T�?�#�B$"A5��xm9ı,N�wzԺ��s&�2].f���bX�%���6��bX�'�g{�m9ı,O~��6��bX�'����ӑ,K����fk^xHKf�%�ŝg�97nG��l�]c#��=Gm̦[�k'���D�B
F"�"��l�\.Y�љ.��f��D�,K��ߵ��"X�%����"X�%����u��1�`�	��<���%�����m9ı,O����h���5I.kY�m9ı,O=�xm9�R:���'u�����Kı>���6��bX�'�g{�m9�?�Ռ"�b�H��E�EL��,O�O��-Ԙj�Ɇ���ӑ,K������ӑ,K��߷ٴ�K�j&�w������Kı=���ND�,K�~����s&����k2�9ĳ�H�!!H Ȏ�}�y�m9ı,N������Kı<����K���,F$b��!Q>����ND�,K�?v~�kRܷ),�Mf�&ӑ,K����]�"X�%����"X�%��s�ݧ"X�%��o�iȖ%�blLGK
�! �� �b)BVb{Ѳ0��>5zL�L�.fb�,�V������U���Wr�X��m&�D�\-�\�ͥL�F�j���:�8��n+���2�.3NzR-P������k�W�x��쵊� Χ�ex�kՍ]��1qVـ֬m0��|�����+e��z�6��!�����d�q��N8ڲ��9�ꙉn73��&6y�G��[�bВ�v�t;2v��ۃ^����E%�6���/���w#>�S��1�f���Jhf6��КGX�������B� Cz�wm�,��55ne�f�ӱ,K������"X�%��s�ݧ"X�%��o�iȖ%�b}���ӑ,K���}�<�j�2��ND�,K��ݻNC� ��@"�,b����2%������r%�bX��~���ӑ,K�����Ӑ�1�R	H15Q,OwzԺ���MXd�$�˴�Kı>���6��bX�'�}���9ı,O=�xm9ı,O{�v�9ı,O����r�uf���Y6��bY�"����1� ����j�9ı,O����iȖ%�b{���iȖ%��)萀�"�# �c�;��M�"X�%����K&��Է+nf�WiȖ%�by�{�iȖ%�b{���iȖ%�b{����r%�bX�}�����Kı;߶[�5��L&3S+��[�@A��''�<�zӆ���ݏ`�������z�,H��&s'9e��S.��Rk0�yı,O�g]�"X�%��o�iȖ%�b{�w���"X�%����"X�%��{mۧ�2f�2VMf]�"X�%��o�i�}�2U,h�cD��B@��2���"�N�����"�$@�b�@�ș���}�kiȖ%�b}���6��bX�'�gݻNE?1@$#AD�w���{���ߧ�+��f������bX�'�g�٭�"X�%����"X��CQ5����ND�,K﻿�iȖ%�bw������L�Rj�ֵ���"X�#�$H�BQaQ=����"X�%���]�"X�%���o�iȖ%��$�O���٭�"X�%��I��u�V�35�K�6��bX�'�gݻND�,K�`���"	�����yı,O����m9ı,O��xm9ı,O������u���cu�)�;]��D;e1�@���q=���]n#��Fܰ�&�Ѻ��Q�����K����nӑ,K�������"X�%�����~� D��5ı>�{�[ND�,Kӿ���1՚��kYv��bX�'����m9?I�SQ5��߿p�r%�bX�k����"X�%��s�ݧ"X�%���K&��&j��s33iȖ%�b}�{�iȖ%�b{���c �/��BB ���������l�B����(��!A�^(͆��6��:Ȓ0�FH0B�06�tj��5\5��`���1cє���F)>ק�{~2���%���w����8�IBqC���2JA@o�a$5�F��}�����iFX��0�}�M��
�'R!@f���/�Ѝ0�,6� H�F�,�S�]4�1��Z���WE}|5�>z;�'���D&F�ҫլbM�M)Vk��|N�������p\�
��>�Y��(�0�|���6�u3>�B`h��5�:̑4���M�q��9S�]�}�i�&���&F�2H�妚�է,��b1���0�$���D�3C�^m|mn��ՠ4<�a�U'b@���3hȁ�M��L���3	�f��tHj���`�TpQ>�=E_TW���b UG@+���
~��:��L����r%�bX��ޙ�_�N2q���0�q�T<���0�r%�g� @�O�����"X�%������Kı=׿w3iȖ%������"X�%��ӷn�N�Y3Y�+�s3iȖ%�b{���m9ı,Ou�{���Kı>����Kı/�}��r%�bX�}��v�h�fx9��ϣ��gt�n�\q�oWn�=Z�(��kh�N����?���+��g�,��Ȗ%�b}���3iȖ%�b}�{�iȖ%�b_~���� �MD�,N�?~�ND�,K��R���L�Rj��fm9ı,O{���r%�bX�߾�m9ı,O����9ı,Ou����rbX�'~'�c�:�	���]a��Kı/�}��r%�bX�}���r%�bX��߻���Kı=�{�iȖ%�by�}u�^����FK��ND�,����nӑ,Kľ}ޙ��Kı=�{�iȖ%��h�	-R��[���]��cFM(F@I ��.�K�o���Kı=�����R���Mff��9ı,K���ND�,S��H_0�~��T��N2q������eȖ%�b}�}۴�Kı?��������M]tal�:�t�����$F�R+0dtL&�0$A�=�7��!�P�fa�O"X�%���߸m9ı,K��w6��bX�'�gݻND�,K���ͧ"X�%����v�u&Ym�3Vk0�r%�bX���m9��j&�X����v��bX�%����m9ı,N����r%�bX�};v��5���V�fӑ,K��s�ݧ"X�%�|�zfӑ,����"dO����6��bX�%����m9ı,Kߧ׹�j[��%�2kY�iȖ%�b^��siȖ%�bw�w�ӑ,K��s��ND�,O�5�����r%�bX���������f���3Ffӑ,KĽ��ͧ"X�%���{v��bX�'{�v�9ı,K���m9ı,H	�F�2b��Q,��ow������mB�\J�װ��t��݆�ێ!�Ց�C�Ls)���ڠ9��0�UU+��>�g�;%p�l����(���|Ż6Wk��0�ٞ�a#p��μ�=H�W<7;g��HP[-j�s�kw؎�=��C�n�e�]Z;9sq�F.ڸv����wCE5�'lz�@.G6��N6�rOR���|ވv6A	lէi\�uo���w�׽���m�ߗ���1rn{#᫰ѝ'b�_E���W���3-�Lՙ�BI����HD��9�:�p��ɓZ��~�bX�'����r%�bX��}۴�Kı/{ӹ��Ț�bX����ͧ"X�%��s�՚�,0̑ˢe�kiȖ%�bw��nӑ�+$#���b_߿�iȖ%�b_߻�6��bX�'u��[ND�� $D"�ș�����/5��f:��Y�̛ND�,K�ٴ�Kı/{�siȖ%�bw]�u��Kı;߷ٴ�Kı=��MɣW�dup���3iȖ%��b$ �D�H�����kiȖ%�b^����r%�bX�����r%�bX����m9ı,O����[�0��n�p��fӑ,KĿ}��ӑ,K�$U���!?~�?M��,KĿ~�~ͧ"X�%�{߻�ND�,K�O�~榿�:�CN{Hslmv�nkr[GqwP��E�Q���cv�z#<Of^6��:[MA�ֳ8�D�,K�����r%�bX����m9ı,K���ڇ��@�SȚ�bX��~�ӑ,KĿ�;f��n[��hɬ̛ND�,K�ޝͧ!T� $i����M4�Gࢰ���G�D�K���fӑ,K�����[ND�,K��}�ND����"���"X����l嚙f���2�m9ı,K����m9ı,O��{��"X�#D�N���M�"X�%��ӿ���Kı;�>�qոe��Z���r%�d��S�� �O���؛�H�w�?�d��eBd�>^l�r%�bX��}�Y��3	�sZ�m9ı,O=��6��bX��A�'����ݧ�,KĽ����r%�c'lnlS/�'8��W�P�L@/�p�ֽ	(맧��o����%�f�l�:s�T�v���=Z�c�י�*ߞ���ŉbw���m9ı,K�w6��bX�'u߻��r%�bX�{��m9ı,O��&��4t���e����Kı/����r%�bX��~�bX�'����9ı,O�>�6��S�G��2����L&5�S�o���X�%��w��iȖ%�by��nӑ,q�H�Z �2&�^����ND�,K���ͧ"X�%����F�b$y���h���_�N2q��34����9ı,K�ӿ�iȖ%�b_�����Kı<�w�iȖ%�b_>�_�\�F��������7���{�������Kı�{���m<�bX�'�����Kı<��w[ND�,K�~�����Ʒ�ۥ����8�ŀnq�Mn�	�^Gi#�Gu
oz���#�\gFvH�33iȖ%�by���bX�'����9ı,O5�����"j%�b_�;�6��bX�'��������2�]k3[ND�,K��{v��bX�'�gݻND�,K������K�q��3b�~s
P2q�t�s��9#�D���ND�,K��]�"X�%�}�}��r%�bX�kﻭ�"X�%��s��ND�,K��K�e.Y��2�&k.ӑ,K �Q5�gfӑ,KĽ�fӑ,K���ݧ"X���Da"�P�6�oq=�w۴�Kı;ӲnMGL���ffӑ,KĿ}�siȖ#��IrB]�����'8��W�����bX�%����ӑ,KĿ}��q��)3�V�Icۧ$�cuR+��77[�9Sϕ��v3;8�jU6�b�Y�ND�,K��{v��bX�'����9ı,K�g�͇�"�Q,G>���/�'8��[��(PtD�$��3Y�iȖ%�by��nӑ,Kľ�}��r%�bX���m9ı,N����r'�	?�"dL�b_�����֥�nY-ђ\˴�Kı/����r%�bX���m9ı,N����r%�bX�w;۴�Kı>�w��p�S,Ԛ�nL��r%�c�	B&�k���m9ı,O�g��iȖ%�by�w�iȖ%�b_{>�m9ı,N���d5ns0�k36��bX�'}���9ı,�������%�bX��ӿ�iȖ%�b_~����Kı1������!�wV�[j��J�Ξ����֍�8'p]g6���;7T�_�mo�U@Tp+�9�UU�뛭ձy�H��d�����z��Jݶ]�8�z� �ڎ�4on�u���s㗛�c8؀�md4kn8�ݝ�ݱ���<�%��qkmmr,m8ӻ]��^�����qx���ꣵfN���[l�&��.z����[��{g�t��uGN�b��+Y$��{3TDNL$A4��g�%�.��t�2uq��Q��vG�����.X�ђ�3��%�bX�w?~�ND�,K���siȖ%�b_~����'�5ı/�~ͧ"X�%������k)r�u��Y3Yv��bX�%����ӑ,Kľ��siȖ%�b^���ӑ,K����nӐ�"� 4;(8�3�PB!r���!ə�_�,KĿw��iȖ%�b^���ӑ,K����nӑ,Kľ�}��r%�bX�k���kZ��&�M�36��bY�D�2�#"g���iȖ%�b}�?��ӑ,K���>��r%�`��O�����"X�%�ߧn����f����36��bX�'�g{v��bX��+����]��,K��]��m9ı,K�{��r%�bX��پ��5��h�jC5��6�kYŹ[�l�o;sI͸HC/��;��F�mJ��6��>{�7���{����~�fӑ,K��_}�m9ı,K���mO��"�Ț�bX�뿿kiȖ%�bw���-�,�˫&�C32m9ı,Ou���Ӑ�C�H ��(U�E>S�DȖ%�;��r%�bX����[ND�,K��ٴ�Kı;ߥ��!�p˙�f�5��Kı/�����Kı<���c��(ș�߷��iȖ%�bw_�kiȖ%�bw��kZ��2�].�6��bX�'����ӑ,K���o�v��bX�'����iȖ%��������ͧ"X�%������k)r�532�e�kiȖ%�b{߷ܻND�,K�}�u��Kı/~����Kı<���bX�{���O������2L�' v��p^}���GO:
q�p�X ���fk�A�G�&���/Ȗ%�b}������bX�%��w6��bX�'����ӑ,K���o�v��bX�'��w�Zֵ2ɬ�D�e���r%�bX��}��r��&�X�����ND�,K����ND�,K�}�u��Kı<�}vh��њ�CR�fӑ,Kľ}��ӑ,K���o�v��c��7HRģ1 FHBB2D�
�	��$a"�Q<��~��bX�%���ͧ"X�%�|>��kZ��d�0Թ���Kı=���]�"X�%�����r%�bX��}��r%�`5^����r%�bX�����r�N�َ������7���{��߻��"X�%��	"��߻�6�D�,K��߳iȖ%�b{���]�"X���?���� �ᔱ�f�)��
��vJ�$v�փ�6���Og��0��M,�.f���ӑ,Kľ���ӑ,Kľ}��ӑ,K���ܻ�	<���%������r%�bX����Vk��d�L̙n�6��bX�%���6��bX�'�}���r%�bX��ﻭ�"X�%�}��ͧ"~��]T�K��ߥ��R�jfe�e�fӑ,K�����ND�,K�}�u��Kı/�����Kı/�w���Kı=��p�;��#5��5�v��bY���RH��������"X�%�{���6��bX�%���6��bX��"(i0@�b}��v��w���{���~�����g�������,K�ﻛND�,K�O� �g߿��i�Kı;���v��bX�'����iȖ%�b{�{rh��MZ\�ޖR���۬z͗^�W�k�-ۮv��^7j�'�·˦���۬5������ŉ|��ͧ"X�%��~�r�9ı,Ou���ӑ,KĽ���ӑ,Kľvw5�KrܲK�j\��r%�FN2���ze�\!�2����7z)9ı,K���ͧ"X�%�|��ͧ"X�%�ߧݜ��5uL.�k!33&ӑ,K��_}�m9ı,K�~�m9���BD�K�~ͧ"X�%��~�M�"X�%�ӿK��j�f\�35���"X�"05]��ٴ�Kı/���6��bX�'�w�ɴ�K��c!!��g{�[ND�,K������i�d��fL�Y�ND�,K��{�ND�,K��߿~�&�Ȗ%�b}������bX�%��w6��bX�'ˋ�촓�X���d���� D���N�AN���"g6�!r�eGd�	t�dB�j	���� H���)��A��B��V�#FLVi,���J:$��e1�מ����oD� � �z@��}��<��ش��q�$��k��!"��9�<_Z@�C!��&��8H�P��4lsr,8g7�[1WEc�9�gf���&�5��g4L�� ��v�7����8������@���2�	q8E���T��6��(kLXI�y5D�����M�__:�_����}rc&ٰ �` I �Igf  ��` m�� T�;sv��9��tg6����9b��5�-�A�<��U=�]g �7H`�!殞Z��^�D�g[�@��g�'����Ku@y���ӗC۩��l�vn��6�G�`�� 8   ��m����l$ l�`�	88  �  $(i���P   oPl [I� l      UUR�#��WA<��+[p�nhB���i`$����s��:i��pc�y�ָv���'�� D���J�'[ؑ���I��s���4�Ys�zU�S�E��^6����v�����d�:5�u�D.z�n���d��ۚ�t���y�Pぅou-��R,\�e�<�v�,�ï:=�2z�j�f��XL����g9�Aɣv�ܭ���ۚyb��[J��,�vX��Dnk=� �&�vtvC��IÃ�)���#�96,ݑ[k�=����U�����^x��N�;3��s�Ijv	�lr�=lnյ��ݗ�Ύrמ�[�����v���$�v�����g:-�S�u̳��Bp��x�\藖9On'�ᛮ9ĄͶ��9��uNj�N������a�8�vȽgѭs�J�U� .��A�$�wd'��[+PNy`���㜑�^9M˺�x;\C���*j�r�n�,M��k;koj�gRm�Ų&��v��6��b�s�$.θv��sؗ���OnzW��Zv{^�{\�S��V�`Oa�طQ�9�I�(kB7ky�9�v�3�\��]q���e����la�ThV��b��΍l�h� G��y]=��s���W��!9S'5ƭ�������8 ���a�n��;#�Ŏ�a��ع��:W���s���n�]H��^K+]��{8P�憺�=��d�E�Z�Q�n���z�Ԥ	�G- \,��p�3���p�зLI=z�1���9z;$��w�����=ݡP=Q}F����� &*��.'qOO | Gh��xpS@�� 
��̲]d3F�+�]�{\n��=@I�z�S<��b@�G�\$M�Hؗ�@.�j���<�n�2�ֳ,�{@\S��5��b����b�9���
�ն��] ��v��4-v-c���J=�"j��[�y�i�^������ƵҖ����u��g��4�<������Y���3ͱ�;6�+�ͻv	���]A#�6P��Ltl�K[��9��۽�Ii�z�-I�Y�N�Y�ς����3v�J�#K�mi�ź�巴���#:�a��w��7���x�߻̛ND�,K�}�u��Kı/{�sa� �Ț�bX�����ND�,K���?\.Fk	5�̛ND�,K�}�u��Kı/{�siȖ%�b_>�siȖ%�b{���6���
��#��,O����u�kS,��4f���f���bX�%����6��bX�%���6��bX�'�w�ɴ�Kı=����r%�bX�v}vkS��3FY�)��fӑ,K?�?�dL����m9ı,N����M�"X�%���w�ӑ,KĿw��ӑ,Kľvw5�Kr�).a�s3iȖ%�b{�{̛ND�,K߾��"X�%�{߻�ND�,K��{�ND�,K�Og׹)*���EmgrS�I��q�o.��Mp�rms��K��;����o���?Wg\<1�32m<�bX�'���ND�,K��w6��bX�%���6��bX�'��y�iȖ%�bt���Du�B�˙�]k�"X�%�{߻�NC�� '(�e���4[Z�#��5��t9�
��T���Y�i0�)p ����B��,N럻��"X�%�����9ı,O~��6��bX�'����k��3$532e���r%�bX�k��[ND�,K��}˴�K� CQ5����"X�%�~���r%�bX�>�e��R��fe�e�kiȖ%�b{��v��bX�'�}�ND�,K��w6��bX�'����ӑ,K��܇�Gn#3$�ֳ.ӑ,K����iȖ%�a�"�c�߻�6�D�,K�w��m9ı,O{��.ӑ,K������Y��J�:�=b1��N}Y�W+�:+�۰�.xv7�3
���g�����{��7���w6i�ᓹ��ؠ/vv_�2C$�@f�R�/�yP��TÓJu.�3@~{̊�&w/vv^��ͥ@��@~W����<X)<jG�[eK@�{w4��~����F�
kS�H R�
�T�q�
�A�	�JRR��qD2���vh|ފ,�w�
"%�$%�]�>fL�=�o�@��@~{̊M��߹ހ��t�re�eK�m 	��Ɉ	&˴7 ?�������3��k1��v��u�f��Tu�U��P�n�ܬ�$3c[Vޔ�x���7b����z�yK��G����~Ͽ~�(�1��8�l��]�* ̼���dW�ɗ$�$��7`\�!|�D �.��}J�2����^�m�- ����l&)����A���	(���-��(̚���2?3;n��/I�(��Ҍsm��=nL@zH���H�5�&m��#b]LJ"^B�&.�NF��.�ѧ�XoWn`�Wf�!5���d���2����i͞���9��H������9��� �{f���@�;R�x�0x��!@z�)Wɛ�&_2d&Jd;�����4m��ұ�Y��I2&� ���&�=$@���_=[>�噒��2�fnN�~�1X#D^�M}�A@z�)P����0u�,QDc�6�rh�t4w�s@���ٹ$�}��b���~B�X���
"��fI�p�2洼��UǴ�xptl�\����:�Wf�y-�����m�j�m�Y�m� =;y�����;3�g �YsCXzS3���cn�w/n@����0�v����^�*mM��ѹJ.:�=�c�;@��aH�Ky��M@uN��f6��s٢3�1�tk�p����^!1qf�n�Mx$c�[�5��ql��eܵE�btd���f�ɛ�. #� C��b�@ DXTT�� @�g���ֈ�fe�Z�A��t��2���5�V�S�5����a뭙ۏ�
f��LL�X�Ԩ��h��O�̗�n� z��C�)�Q
^$��@w�_3$�a�əD�t��������QLC�+M���&�=� C���րw9��p��-�Z�).�5�d�R�C32Q���P�Ԩ޼���;�>�h�	�clx�'����h�n��&d$&2Bd	������t�=����F)���1��\�1v�/�]��5ʏ6Ջ]��]�j���L�#�D�� �;f�{�f��-��9�����ib��1�̃rh���o�Gj�bipQ�)�BL$33��7w�P��h]�K\X���$M���;m�h�n�5rd2HI d2L	4A��4{�4u�Q���� H�F����h�5 yɨ	�+��K���j�B�I1*�3ד@jnC0��	0��J/{������(�%���d��:"��������Ln��a]%Nmn'W��^��9#�N5�z�r�N�crE�~�M ���ye>��w�}r�ڣ�9��1�4��oي?��`�X�bH�d�������������h�Be���LO�9�&��d�@g����R�Đ�3�)#<PaZ��P�~ �EL23	��ɠ��hX�!�
�ɗ���$���O�9�@��@�I��y�����*�iLQ2H=feܒy��f䟐�X��H�b�^�<�Ξ(�^=�2a���<��;��Q�OO���>�[���a*�� t�8y-��x�Dn�VZ��:~�z���r�t��s
v"J���(y����¿�ə}�L�0�0&�3	L���= n��4�ڦ�{�V��d� <Q�n�/�=�ɣ[����$0�HL0���s������J��Ĩ���Vf�� �P����A�W����� ����s�}��s�r��$�1�!�4�ڦ���p�2��������fM�}��c[���-7S��[Y�øycؑ�W��Gz��v]֭��\�x�x`�/�c�M@>�- F��*����������l�L����<D�~�ǭfe�|$�C!2M2w}4���4��7���H�v���(���R9�}o�@zܗ�t��}�Z��.�m�˖��֦k3r~Q�`"�":�7��;;���E��]���+q�T<�&�x��d�&d˓$�L3a�d�d$�������M��0~m�����z8w)(D�a�ۘi� a˂�v�z-ӝ���<9�mQ/��3�5UT����9�����.��H�s��^�#U��6t�]v���ܶ\�˲)˩��p8"qP��BtuR�y0�a����<�3w�	Qđq��:�=n�ۇ�a�n1�n�/9�t��H�.s��Zv�sюM��.��K��.ݫ�0�'K�É����~�~����i�74\�ulk�o^�q�hT݁'7[�s麸�[�,m�6N��eU�Vɷ�w���- F�=nK�:M@{ΓQ9��S&ܑh�l��<����$	�b�d����������w��h�ܺ�6I1�x)�)&�����O�<��w�[��.��QByO	����x��fe�L2�&��
#��h��z ˼���S�;��o�o��InM��Ƞ>L��3g����@�ɠ?\/�G=�5ڍ����Qڥs47g.��(�l���k2䴄����		�s֑�� d�&����4+ڝ g�'�̿8]���Y�;�K������<���Ǌ���'d�2H=�4�^= e�M|̒_3$33!$��7 Z�!t�� �e���;�K@����� ���fffѹ$њ-�]��/�	��Pa g{������w�z3���$��LK7`��@���@��jz�h�h��U�A�a��#[��َ۱��kϊNm�Fʎ:�r�;�Gh��{��{ �����MpٽsWZ���4K�1� ��'�^;V��;V�W{^�۝	�x�LMH܉��ՠ{ј�=�E�Ǌ�\�0�L0ɐ��Ӣ�=3�/3#�K�����ks���5��0`&�t�B��F�@�
}MH������q����bH���<ʰ�Ca���
l�H$I��`Đ� H$H�y��J%�\GƘF3ٷĉ=���=��x��l�4xL��v	7��$k�>���MRƆ��6o@]$�it�iIZ��`i�	��$�FE�M�K)��<|л���3MT�F��M�DZ�"p^|��
)�5�.	�0���SA]:���!+#	��� ��,a
0�h�� $ill$ ��:aFd.ʵ�c3��n��p8�!g�z�h6Q0�'��iB.��L
*X�B��> ���Q1���z�-G@|��R��_U��Q7�_�����hw�E��$�q$�t켚��(�N���	������@�}�𖸱E�H��ɠu����2�������y4����|��������b)�$��{x�;cr�wn��\���΂�w-`ݻq��ηF��8�mX��^<�O�/"�.�'��a�f�5�y�,��
""% B��p�8�k���3o�@�ߓ�=�S@�� �bX�H8�����<Q�/��2b"�������]��Zl�9�1I�uw�=��M�<�{��"�`4Z!�!m�߳`v�	����145�@��S@��0�d�3=� �ޚ����7��2
��)c��ۭ��tS��Pr��+��X�F�Z��\�g�u����j-ۻ��5 ssPc��9�@Uޱ"��n NM �{f��<��fCDѽ1@^��@�ɠ?,�s\X��dR&�rh��=��M?��<�#�~��~�8̨��(dJjM\����"#�@�Q�9���?��~��4��+�@=8��q(!L<�ʠ�ɠ>Lɒ^l��3f(޼�@P�́3&�2Hh%X� �~�%�Z��>5mԃ�}M]')d�!�^$�o9�����e��0k��YА��]�n[s� ��gn�-���y�n��[�,vz��v��L�.�t��'Wi��X�>͌ �-���͈�;U�Ӄd:���:|�_i�J���̧.{-�N=E��������m��Y:P<x�T�:��q��s��tκĜ���k��h@g�x�=5���绿������?�7?�2�.kGe�G��sv�7Ql�z�_\М\�kkD�l��%֍h3��,�3=�z<�s�5 ��rt����9_rb����_37�s6h��b�"	��P������ɊԒN�6� nn� ~���̙|�`L�$�A{�+��Jbhj������ ��h����Ǡ\�.,17�1�$Q��o2h��&���y1Aɓr�Ɇ�����?/�b?D@�2�
I��hq����H95�������[j�%�ĖzÓt�v�˚�6G�����;'ZU巴�u���e��o���&h޼�@y��I�ɛ�! a$!��W!���P�/�D/��K�����?z�gɒB�(�vh?o�@�^�4Ӂkm�0s��R* ˼����(�K�d�C$!$����7��@~��B�%;�"b^G�����\su�qR ��@wgn�4�q�xԆ'#�8�l��fy�$��2l��Հ}����ב@���.��T+q���)�7lG7on�����bS\7]�.��+�;.�N�pBm�n�=�*@��_9�����X;�?n��jOMK���D� ˼���/��C$�D��?oL���*-���$��!I4x�Z홹�kCj�� �*)ҁ @�)"��U���}ݛ�N}�f�rڍqb�!�H�Qš�<�<��0I2Q���4f�* ˼���1�q�Q���&4��h�n�^�4x�Z��ɠg�y���|4L�Da�u���-��X�Z�
n�Lgj�Jd����=GmԱ����y��o��k1'0���ɝ ����h\��W�M��s@�� �bX��)��@9�ɠ<�y3@{ٔ�.�kY2\0��aB@WZ�|~������f��4�&��_��&��[����@9�f���&\ccn)�$�C�3�<��{�� nf� {ٓA���Jf������3H:X: hY"4,�A�)8�L	��H���5�lJ�B��A��{�s7$���mԉy����@���̛�2a0̐$��3;��k����fR�?x �&`OY'u��l�ۥ�ȇ�S���8��s��Iջk�87&"I�"JI4
���^L���_3~p.�f�՚k�����&faC��o�ɚ��!0��C&0����Qgu* �ޚ�"��Ď��b�ر�<ۀ^[���\?��<Ī�k�8��I��:��<&�̹������ @ D$4Fn�����ד4{2���H�bXڊ)�I&�W{^����4�e* ��M�&^3�:@�$�ݍ�������\��*հF9���j�m=.鸎��mt��� �n��&P.�j����N<�j��!�O7' \f8������r�8.L�ms�K%v��ɀϋ�S�^];�m6��\ڷ�;6��u!��K�[�*$�PZ�ݖ:v2=��Dɵpp�ܾy��0��OM�U�MuC]��qt����.�q�f9;YY�sWgB'����3�7f^}�s���ӹ���ӏW,7Z���8�ۚa53)���N��,H��"D"�v��w�?���7L�ݷ����n�'H� ssPۘ��jV�n)��$�@��s@9�٠U�נqs�M�ކ\�����I#�]���y|��ɗ�d��3!0��	�$�3�������E�)�� �q	�4?��_;~zWo�hrנ�l�.s�M�kQ�ɍH��s�~��'��2,H�"�3������@c��P�0��$8<ʻ)"A����v9^}9�5�V�WS�<Sn9q��ڑ1��8F8C	��h�ՠu��({���~p={�4�Cb%;�,�3Z�]�=�����U�q�M���H����Mn~�w�� ��ߔ�*�@�� <���jF��9�W{^�{�T���ľ]��Uo�@��P6�NcƜ��C��?y�g�	��BL���3���4Ͽ}��������2�qD�9@K�1 �	m�@�/P��������M�b.*��I�v�O�]��r�����E�d��t=�.�wy�MC4��E�y�@����I$�M��2	�$��$���������b�p7NG�U�^�{�T�*�@��k��31#�|&�5���I䨘��^���y�G�d��(vt��H�L��Ij��B�Uټ�M�dF)P�@(B�+��ˆ����S�?�� 	L�&@�ɲ)�>�_��(d
���1�L`�S@���W{^�Wmz�-S@=)Q[����jzɹ'��~����~W��E�1�0`0��b�����k�'׿��[��h��ffs�kdmō�"�x&�m�ׇ����+d���y�8�Tۍ����9c�d`�
bM��(�~��|�W-O@���W{^��W�P�ND�<jcw����1�3$��nl�@��@c����T��AD�##��302L�2o���DK���������7� nj[��r� ����1���) �;f�Wm{$��߮�'}Q4�O��#03$����P��AҞ\�B�"\y���& =m��s`�;���S�d��s�6tGVz;����tJ�s�/���3X�Ȉ��modyuei8K�mf�����9�@�j[��3���1�a�D��)���b���%��@s�tP��(ҔJ�1)�5�R�v��̊?��'>f�P�:P�d�,S�C�y������Bf#�{�������h9�4gU	4�NcƦe�n =m��s`�#sPܘ�c�HF)�X$�0�#HKB#u7�H�%aV6d���։H��[$�.���D)�� a���\�=N1��$bDO#�=����� hc�!0`I#�JGqB$�Á��Cp<H1!].�$3^H�p"{�� ���]@�6��/��g���t�
��1߰>HSU��ױj`ohk`SB�=
i��AO|�О��0	x��^��������G��l�̅U�P�` H��{\28Z�ж� �  a��rE�d�A�v��ΗN&N�Y6'5Ƿ`��p]f�ێ��{<\��j�CڝC�<�1�#��[fP2��}�ӽ��S�W��i�0p�kC�=��c��7M�y괾��� 8 � -�m� �llm�[@[�p  �  $
P�$�v    ��� ԁm�h       ��i�]w6ڥ���=N^�=�n�����'�p�.n�khu�`�6�ӎ۴G5�Rv��v���fS�x"�G���sU��"�i��g���M����i�rp�'(��%h���qz�%���:\��y�ti) ���ܣ��N��:xZ�t�3������,�;�60qgq��Q��褡�`;�OXA"��ܵ�ȝ���:�]�P:h�]-R�jK�dKdN���4�Zt�k�#��δ��$͋E�����vv�;.=6�[cgL�v]�j�H� ��mCŭ��]�#n�$�ӈ�K<�;�3�J̽Oo]��:wE˥�N������u���f�m���v��5�6(;u<9r۲\���#s�pu`�V�ӵѮ��.��4X��x뭮�@��L79�H�F��ۮy�ۊ�@�$��({�0D�*���pЫ.��:�NY{)ۻfثFkX��$7����������m��*�ng�8�:��6��4$Rm��7��(N���:�q�U�d����l���a\�Ӻ��kg�ː��K�r�g�,Γp�F�l�&�3xx�+�[��L&����c���L�]���Dn)Xw͋�`��7f��\�����1����ć<�m���ڶ�c�ݚ�r��x������й���)<<�;H=v�t��\I� ���V��h:�f�gW*�Qzg$����Nv���'[�8yx����]m�:\W[ON6y�ĉ;�۷��=N0��d�3���3�������'ȬA"��g�pbbЂ�T~UW�C�s��fM[�j8 *㴩!���>��v+��㗴gт�gf�¦v�j�ٻJ� � �UR�B�rp��&ˢh�uc
7K�NIW]�o;k��ݳÈ䧇,�.U���痘
+��������an\Q�]��nL���K�5�Cu!29��Sr�\���N��r:K�E�˹����vݹ�����7�s=]n�=�����vd֬�j�S2g1T}MsvKy���7;KM���q��ܑ��c���^��d�^7a�oQ�&;\�����m��N�y4=�F�@̑�}�x�>Ͼ���1�#�R{�4
�k�*�jz����<�>���LQa�n RM�~��w�=?g�a�Hf����;w���3���O)	<��@�����S@/{f�Wmz8̨��1�a�D��(�����& %�/ʷ����К���I͈�����m��S��V�9v麸�[�!	�g�g��f�=4K��% �ic�@�_�=���
�ڟ�y�fg�>�O����
bM��L�{$����ބ�
i�`6ƅKk	
�D0V+�K>���$��s�ǻȯ��@&DA�#��"e�T(y�@����z�S@���@���u��I8�~)$�=�)�c��P���&O�����Z�Q.�yrb`y��ǻȠ>M�cz���r�����S@�w:2��hLra"-Ǚ�Gj�:8hn�Vx����J��5��Z;#�F2LQa�n,�@�v�����v�M�����m�kS��2�=�<W7	$4A���ϻ�@^Fc��ɝ˸���`�%
T"&^(ݝ({��5%�L�Hd������
��4���s�rNߏ����:%[���F��9��Ͽ|�͝({W�A����f�f���|P����LI51ə#�@�l��Ws���S@�����~7��x�%���n�pvu۲����觮�Ѱ��K'[�ש�a"�r)1�S ۋ�>V����l�@c�d|�|&a/@f�����:91$����D�{e7�<�>W���@����-��2��$�=�E�ǣRffN����@{6t�/_X�1D9�1��N=����}��@s����2p�t�2����iLɲg�y����j���Q�i�$�P��x�>L�۵��5�v(��z��}/�=��_6`Y�NBx��v����n��F���AO)�`ݬs��ηF�m9�\Lc�?@��O����������Ì?+�����K�sq(�X�!�U�1 �Ih	|���� =��ʅ�I��&d�=�v��v��߼���Dgt�@s�tP^�s��^eB��-9�W;S�9l��Wmz�ff+g�-��,>�$�Q��H���eܘ�o$��9���aﮮ�� H��d
z�GA�H�Hh�4[ I$H��I#F�%����<��f�֡�;���U��YZ���q��6{nx6�6�x�s�T�_�mo�U@VҼ�3�5UTvZJ$��^xƗ��v�4�uS����ፌ�2@\jgVnݻa�ꮞ!���oXWHY[���-�
�cmyӭs�]��N�l��v��Z;h6���޸mr(t^nnF2����=v:��ݢ^v��2�ۮ�&��j���t�l8�t�WE��d��
���3f�j�TIkV��e;Te+Jp���q��{ւ�c��^�ϣ��w{���۾;��닝F������䖀��7&�[�LPI�!�łq��h����e4
�k��<Ď}O�{���O$y�z���'
>M�̑Ͻ�@_���@��ʏci�R-���|� 9䖀��- x�s3j�	yxwPD�@[��(n�6���w����=��=�i��M�%�c��2�/F���tַg�z��iN�:t�.7\#�u&��
bM�)3$����Z�����M���@�rĨ&�RcƤ1�eܓ�k߮�Q�"�̒���X�|j�:H5� � � �Э�
&�,]�``�H j%D��T�I�G�}���|����_$�	�
 ��q��t≘��E�w���us����v��Z>w�{r����d��"Hh�s�K@zc���6�0�m<��(gxt<LPq��̾3!_V�\��?W;^��W\oŊF�E݂��9ó��]/o�cdm@���O	nү$i�!E1�ӆI"�=��h�S@��k�/_j�=��ӆ<���ݴ�@;�19hLr���L	2�0�ߢ%<Ļ�@∙(|ފ./�C�`I'I�!��R�@"�(�F�|ڎۮ�h�e4����bI��L�$�̙��rs^���k��(^E�t��jE&<i�cqh�)�~ϐ�&Cvw�<��E��@|�������MԼ��n=qO��C��:�z�qӲ\���6���s��f�v��1�bd��Δ��E���3&_�=�:P�\�L��e<̔��EyjK�_	�2U?|�}��P�@�w�;1A,sk��;��Z��h�S@��k�=�v��QF�OJ�ʹ�Ih�� �*��}���Q�(�'��߷��w$���Fk�5��&!5"�/]�@9�f�z�Z8�Z�gzB�<S0I����n��-�]֧aF&3�9]qB6\����.;z�g�(�����女z�Z8�Z�h�ي�1$��&G$���5�/�A��@v�s���4��]\M8)1�NbjI�s�ՠ^�V�s�� �h�X\bI�25#��.�1��̚ �fMs(̮�;�? ���Bx�19�s�� �h�h�h�۲&�p���W�
�E�&�)�7%O7�L#��⻴�HH�j�d�m�]�n[k�`YbY��$G2���afh��Wv���9���s�/Y��(�u��������K[�m��]�ȐY�덨\i�;��ȷF�#N���ݏnq�kc�qGu�j�/5�Hܽ��5��<�r�kl�"oF䰽}]��5�t�w�/�[�Y��&�h�=�{�����ttbjӝ5|�P2��i��"v4����0�I�ۯg20�W(%�a�M�8y��@��@�]�@9�f��s���ģ��i����=��z��(�v;��3;��=��_�M��ߙ��y1	��k���@9{f��;V�p�TiW1���qŠ�@9{f��;V��|���b�`9�&���9&�r���$���t��nn0�sh�yy�;�Gg���܎0/D!�ˣ��`M/N��:ciۗ�˵dX+�F�-|�?�ߢ�Ih�&��j�K.��]޳5]fk3Yw$��}��)1Oja�)��cKRfIj_*{�4��4��_32L�^�pZ��\xPLJ������@�s� d����0��hNI���@�;)�_�1�9|��@^��x�gy�QD�����̛.w_��vh�y4�ؾ�m��O���i��Jdn^�����y������F]����I���F�mqj�ڲ�sO~�h�&��j��h%F�sd�<�Z�-����@goM���~�ǯ��&w6�J���j8�E$�߯�@�;)�λsF��3�!*k7f�3�ˡ1���)���Z��Gӈx�	C�I���� G��A��ִ��,=f��,��8��������9�p�����5�\+;>)�5`B���y�S!�C5�֊a��SF��0,�R�Sf��
��ˣy�1��ύf�����i��vl�HMBN�v�th.�U�
p�!�<a��jh}�0�W��u�OT8i�1'��57���3Jߦ������#�ĸSFzq�����<�S�֭��|8OI�p�z�u��8��j�rm���0�4� D~W�਼ �_<}D�"E�!�L�� 
}O���C�>TCB6������[UK諭���l� 㚀����JLmH!�4s��x�Z�-�3|���@gG8뜇w"f�f	��K@rj ��9���_}U�?�w�}����e��6"鋮��&���_S�s��r�N[v�'2s<�ݞM���a����~ �����j�� d���^�,���Ě�h/l����"ݞ(��z �y�@~�o�L�1)�Ӄ�I�s���;�j�{l�^٠s��1	ىCLB��@���?^d���h%&Iy7%�Tn�� ��|��M�i� �qh��h�g���_��v��w�ՠ^gc��qck�9�slk�u��v�)�)e�4�z�t�sWn�q��x�<Wl�L]_6����5���K@rj�v��/2�%93@z�p�d�7�4��|�M ��+�ex4��k�#7t@>�- yɨ������P\�$Bx�jb�- ��� ����
Is2#r�����!)�wQ'�ye���j�� d��<�ٹ"�$�ʁ6�B(��
؉*��@�~}���s.kZѭf����n,/<I�۩��
T�c���R�EƩ��W�(p�� �US�tc����D=a�3�-+r��+WOOb}�7��^��μ�6��ÎZ՞2�K�n�i�����M�Ξݓn� �{Ԝ.�6����>�m���#��An�c�ɶɭr�x_gugM��/���x�q��t��K�=qv��y;05!�uk{<4�fz�lQGw�r�Z�SRh��5��GN鸔����_3�㮢{�y��Z99ں��{#�ƲG1$�D,�7' ��|h� 95 t�P0eM�Jͳ���䖀<���M@s{�*�4@Y����"T<�
&%���h������K@N��sh3j�ڎ)�I&�r�4w��z�Z�m�{�AtI��s�;�J���/�1����3��hٙ4����m�x(�Ǳq��:�gݺ̅�_[�c�u�Z^�d�u.{��oQ�!��1�'�t��_�- ��� �}��y���>4}�b�|�'�6�)"�{l٘� H��"�Bl��iI�M@_�ɠ=w8Pq���s7ɘ�1�]	���;����ǈ���呂�w8Q�L�;�F���6h֭�fX�(��F������\�~4_�- ���@9m��N�1�LP���@��Ǡ9/�����wt���
�����m������bNdc]�u�^�n��<l]]n5Ϧ��z���cd�h�anGV�nw6����:I�7��W�W�$�߭�s���$��)�G&�r����<w=�:Pq����&�&o�Q�k������DD�4n��3�fj�`J��hJ�� �W�4��+�ex4,r5㑎G��L�s���ݚ �^M��y9��;�}�>��D�%1I�{�f�{/&�������zS$ͻ&l9�rƣk,m�n�u:{C��kTpW:�OGgWyn�9��p����???.-�ͼ	�� ߻�=qx��3�L���ݚ�*�\���1D(H��:�V��f$^��Z���@9{f�s�V7bA�x��h�h��i��g�e���_�ߖ�p���Ssd�0�Z�m� �^M�Ǡ��fB`�I:fY��%�@��ت��1$�qL�I4����Z�Ih�M@z�6_K9�v�d���f8:,n�zΝ�!������٥�����u�绿��_����쫇����}��w�ՠ�٠��@��R�A��&�q��zx�Z�PG5��b�O��/�n���h��@�5 tsP|� d���Z�Y��8x�BrM߱����@���@_�1�>I�w�����aED��(�	�@��k�;�j�yl�^٠y�y�[J�I�ڍ���F���9�<�ԍ^-����#T�'4�ae���Z�H+<HR� � �UR�\� "w.�����]�V놜�ʵ��^c��#=r�v;R��^څcbd���3]�6�׊�a����H�#�[7]۸�#ZJk�����M���G/�g]�:���6'��F���n*ʒ"�u�z�M�H/f��e-uX���ֺ�8����̽=�M|1|فg	r�ǎ #�3�Y��d[����mU�:.,s���h��F:�lc��}_��@=�@9{g���aU���
_���ɍ9��&��yl��j�������ڲ���Q�2)$�^٠qs���h��h�uD��)!$`7&���ؠ/ј��ٓAː�3����Q���KMx�n8��ڴ�[4��h\�z9�$v�M6�q��&t��ͯ)���γC����kA:�1���+��ǎy<�'�Ls	"�yl�^٠qs����=V�Vb�%��؜�I'�{�o�H���Q�,�q6*- C��~$ �f-�^���~4�[4������!BE$�8�����i���G;��@/���uݘ��b������̚ ����HI�f��ފ �_5��y�`�4�[4��h��Zoe4y�`�p�"c���/F���ttϭ�q�l>��6�Ӻ�;����y�Ĕ�!�Ȝ�@;{f��>ՠv�S���\�Ψ����$$��hz,�=~�(=�4yy5�K�|�2�7�;�� O��/@w�?I9��f�B,$�Zb k���=��Z._\�$I�DLnC@?{2h��hz/��I�7+J ���pı�Ě�hol�?��?�����~�~4�[4w��7�Q8�݂�û<�L�o�"�*^�m[��k�"�qx4�D(BI4q�����M@9��vVdڲ�L��2�e��d��٠�٠=��ZÆ�SD�`�4�[42�hԒI|�̦wc�z�~(��$�	H�D�ol�9�ڴ��Ϧ���"����PP��ĀD�T^g|��t��~&�ؤ�I�$�=��h��h\�z�v��:�Y�̑�m���/"�5J}A�\c\�z{sb�NУ<��v�A��-���׎7#�@��S@���@;����Ʉ���@g-g\��]�;��&D�s�5;��� 4U%�$�NG��������hs���U���OB�$�A�������������P|�&N��呂w������sƔ�@�� %�$�P��@]W������BC#U��1�T!�c&� �w�����Z55�8B�H��]`����$hj f��h�X��ӽ	��فZbA���B$!RE�# D�)\���� I�u`)6AVҸkDE&�tB��"֎���^BExk|%�Vc�'0v�k&�]h����
D B E",dA ��$����H�$
�
�R Oov����{����]���c-TN �` H�R�V� -��m�    Md��A�b��P�=�ti^�.$2H���ӭ��c����9>�v��i��y�9����,	���|���o'\��AV�N��ɘܸ흩Ҁ�%��)�h_��J����ز  �  �$sl� �c�-�,��lꚜ   �  �)@K(�F�  � ��  im$�        �afݥE���c _2�7;�٣lU�j����Wdv�w6�c։$vy��v�ym�kҧ��m�f�2<i�X a!����:cc]Hk�+��C�%�z&��YZu�ע��/W;\�c�]���������(�v�1+[g��=��g�������� 鸱��� �7Ϝ���,��r�ݍL�]lk��r��X��bܚ��{*�θ{#�9�� YV50��N����N�n������۞D{��-�8���#���<h-=e]*kp�rqn`]`����3�����闩V�2��hz�E��b��9�B9Ӧ�rX&e�eX�Q���)�lix.-fycCU��@;iP��n��zXV�n�uѮi�V��vd�^��"�*�db6p�����$�J�Wi�I]�� �û'�v��Aw��0bһX����L�73=�:�B��ц ��(�Ix���1l[��M��*�N�ufAq�� �=�.������6���˱�Ά�%8���U��v���3����g֩��������p����l;�y��m�{��צ^[��+6�њ��d�ۋ��#,�M�[P%9�tn�M�̶wm�]N޶F�s�����u����ero�:�m	�e��tѴ�x6z;X�����L���R��c' �nv�*��)�n��ny��q�2�[m�� ��JƎ��.���WG=px�V����n9�p��6X{[�.a2���>�$`*z�A1�h�M��(�SB x����R�� x
��	����`v�＀�U�m���Da��ې!���� 5�T�Vh۠*��'t+�@gY@�l�v]��:���FN�NZvz��z5���ڼ����|������E�z�f�f��;$'AZx&yLA��1����m<�@���3�q�ʼq�8�d{f���Aw4�����.�J�q�/m�C�ه�-/e��mܽ�nc�ڷ���Fvzt�浖�	�fa�	�d�AW�T<�������������0�����K�j�ǣ����:�N�gnY�oZs�b�㑼����m�@�}�@��h������$9"y#�h����c!���z��� �^M�V�lRH�ōI4�ڴl��^v� �٠[����18����qh��@�ɠ�ɠ�䆎��z�s:�M2�	�`�2Pz�h�32g�ݞ��]�h�M�2�12a�'u�)����*m�/cA(�i�x����Ӷ쌩�"��j'#�m�\�E����ɗ�{͊צ��K�(�G&�W;^�y�E�S@�s��fd֦Is|�3)�ߗ9��HD��#�?����U�נ���v��0H��cNx	�@���@-�hw���M�U�ILq<Q���f�s���)�qrנs�1�B9���x����X<C2;��l \����u�:Ƙ$� G$G<o�}�3���t~��c�E&,jI�~�{e4.Z��٠[����18��ȉ$��_I����;������:g�,�7�x�dmHh]����'��Z�it:$��H1!$ 1 23SZM-Z�B@�-�m��u4B$#4���<�����gf���M ��Z.(A,�����f(9|���� ��/'
�����������P�rh9rh��&̝����� {3&��FA�]�X{a��t�
��gsy�������n��,�xЪs�te�q���wEMw�@y����:���B�w呂���_'N��X�%�?�"�/m��[4�j�9�uW1%0HjA�G��� �-�z�Z-zhv��c�E&,�@9�f�}���I��ﵹ6 �*cP �WM���I�%@�H#(��i�%�B
QKD�H�X�*��>+�{�����}�%��f'^9$��h\���@9�f�zs��51�7���^�]u�bBݧ�u\�q�]��]m��������?L�H�B������^�r�4��h�h�z4\P�d���NG��� �-�z�Z-{�~1���������!Bɠ��4��=2d�o{�@��@�n<d��H9�fE$��٠qrנ�� �-�W�.,Xә�4ܚ-z�̚ ��&�.�&��d�&2a7n�m����{����}�X�yW�U�`�,����ι��k��^c�&w(���H�Q��ey��e����6���*��s���6����N�s՛�89ힳ�͸�;�ry�%�61ۮѫ�Ż�d����ˢ���ɞ�D�'5m�xX��l�*�j�+���mv���ƒ��e�6�תr�Jiʉ4�i�mX�2^��t	r*�l�<H]����걮l�o�|��ϝ<ݭ��ꤘ�:ӛ��6Ƽ&�;��7K�9�uKgu�Cn6�ړs��������"l�����_�~��[4��&I�~p��ؠ3C$�C�A3/2�C�� {ٓZ�L��37f���ؠfd�-�R�A��My$	$��٠qrנ�� �-����˛�4(���L�s'��ؠ�٠{2h93:�呂p�h�0�&!7��-�@��1w�}= �女��^���*�NCs�.e��t�J9�����|�b-�V�yu\q�kc���E���y��G�ŭU� ��ڀI���G5�)��u!��K�� _�&���2a�ѡh�
?������rI�~�nI9�f��ӧ�ˋ4�a�7&���^�{/&��$�;�{�@{�@{я�)%2&Ȧ(���٠�@;�f��]}��_��?�iI���&�=�ɠ93>f����b�=��@{��o�@�G��m-Nm���n��nG�u�!{��r��`N�j��7O�kp�����n���_I������1�r����"M#�M��� �h{�� �̚�fnQ��ry*e8��3��4��"�fd�320XdP�v�$Wj����}��ܓ��~���߮�o1x4�D(B94.Z���h\���@��'c@s�)�e�M�2d�{���vh?�"�Ի�߿{������|�\1#8c)�c���<T�o`���k��l�]A�l1�w���|��|�F�1�����M ��h\��Vנs���2&Ɋ"(��@-�h\��[^�s���:�:4�$�LL�@��@�����h�٠[����18��8G������?��E fwM ~�ɠ�J7��3��p��b��.��ϵ�'�4�ۙn�6�M��@�j ��P}& �~�;�(Ϙ�И�mAr	%��Q���
�mE<α�tvuq�-��	�ϓ�VMqn�$�&�$��s���8����v� ����ڞ=�x4�D(F��;^�H�����M ������'chf�i{��w�b �I������k�=])��ō9�xۏ@=�@;�f���נq[^��:�ʔț"2dQ�&�w��@��k�=Vנ�٠s=����䲸4�&�x�A�q�D)�ݻ�llW.�Ѩb5�[5n974�T��W�B� 5UT����8�N�{l:��޴U��:˺���8ἛvGU*#�y�h\���m�A��Ӭv6�����G���y��k�,����=X���ld���q�s��d�^[&�.�%�rn�M���j�)gk��'!{m�� +��ۅ���\rfS2(	�OЈ�oɞkF�5ri��i�[r�N�����	*��#�.3F'�6./O;�,͐�Q\:�������@z䘀=�j ����up0�q5�p$�@�v׿ؐs�}4��4?�"��I'sqc>�g���ĩ����j ��:��@zܘ�<6e�0�&!6)$���vߦ�λ��=]����;jx�E����r =��:ܘ�=�j �&�w����φ����8K�,;�t ���������9]�j�u*,������N6�ns�����~4{��o4��h~�|�I12�<L� ~����,L����Rd������4fm*��@s��<�L��#&E�h;l�=�n��%���h;~�yUf�'#�2�LL�k$̟כ�P�:P�^M w���Kbq��RL�9�8P���6 fn��ٔ�� ���"*�����W���y�<׷L�uT뮠�=%������RF뛆� ��������`�<F4\P�d���$�@;�f��m��9�)��l�9�W�\���������2���f%�gL�lА��R�R
��"m�H �FA�*D��r;dQ�bP'��8� ��6��8,.;$VB�B+��ڑ��P$5����I]o�����D�;� /�X:������FyC�h�+��~i��R0ρ�M`b$؆X$b�Ԥ0�p��3�i7�j���:8�!�DЧ���Ӧj��{.��>��HE�Z�h��� D0)7j���w � ����K���Xl]|n��0]a!�.� BNkI R�0Jiܗ��4���}��D��#H3�P�&��T��d��OC��x2��w�&����D�0T~��>� b��X
��@�����`:C�t��C�����3rI�{�ܓ�����c���$���o����ɨ9 <�S��sv����@��$���RL��~�����tvX�z�]�=3�Ds��u�F��v�"�t�e��L�zm��JI4�f��m��-v���z��M�"}$�qL��H��=��-v� �{f�[�4�u,T��2�wssD��nj ��@y͆���|W7�Q���- �{f�\�����@2�ȶH$0��2d� H!�}DS�x��{�o˹���.(a2LBl�I����y�������뼚�$��_D�8���v�QÍ��9<����\;��o�����k/3q��f�ͷ����@fE����u$��w6h5c�q� ��&�H�Z�V�s��@3/&��y8V�L�w/#F>&&@��z �͚ ̼�9$���:P�~Z8�<�<��#'�E$�ol�<��#� njq,�l���Ȥ�G&��l��k�h;�4�f��y�fd�^$T�2�LmF�JIwZ���)lۮ�dp����וi0k��m (�������������0V�d��.�vWNi���L���v���<�i]�'cT���q�㙍lK�s۷V촇+m��Β�j`vs�Z��s'oD�h�!Xd�^�ͭ:sͳX�</E�����t��u���_�=�.��Cs������u�d���q;���*%n�uSy]D�^�]�<�8��,����<K�Mg�8���y���<�n� z�&�33'��z����^��_f���E�- �{f�[l�=��-v����|�h��"T�q�31@��@e��F�,K��-�~���^=s�OB�"&h��(��z ��M32N�������A1�Mb��@�ڴ���$�Ps`����>
��6[
�Vƞ�e�ǣÞ���'oO ����
3�b�I��;�4�٠{�)�<�����;�G�$�'��\����O���ތ���@�V�T%
���� ���禁��~z��4Τ��$��'0�S13@_�p�1�2(��egoM ~���^�b��N!��R8hv�@���}6���%/�.DH��@9{f�^�4��hvנ{��e��28�#?� 0�%������g@\�����&ǣ��g&TD׋v�LI�I&�^�4��hmy�z����}~_<z�/�(��7&��M�U�1 tsPnj r�������G4��� ��L��A $! ��Pҋ�x�@7���٠w���/,g��^<�,0&5#�e��^d��x��̓�݊��<�'�<y2`E�h�@�~���b�|���h�1�d�$#�{Hs���Ӹ_cK��e�-qα�Q�ݻt�c�#�� &��4�v^��m��_���	V�� 㚀#�P�K����C1H��hm{�33�H/��\٠/"��RI�;����I�&\�y��Pnl�^dѫ�7�y�O�Ѡ�u4\DXL�h�I����/�����&�IВq&��ͩ�!�z������;�o����4̸^�u����s��rb q�@�4���l�x	̃&4�����>���m%vk<�1����wH'=GC3�2`ԊE�\]��ol��f���V�yc<*��a�1��v��95 �9h	V���B�]�LM�Ʉ"�M ��h��hmz��4
����@�q9�y#�CS33>l���v(��h5��w�ݚ��b�1��3���qvנ9�95 �9hV��Uu�����c�%P*�u�]�O]�ްR-ٺ����٪n���m������o�'� ���K��v�tNf�'Y��#֛��J9�b�Z�lv:�N�\F1��CcoC
l�٬�v"����:��^�{�hV����ԑ��˹q[X�c��mΝX�<��z��j[uc]�]nv{v{v��y�ݵ��˶�y��+�iŮh���8��w�����s�z5v&�ٱL]u�b��T����h
�1�Cɻe�����DɈqB(C"���呂G&��-*ܘ�=��,�f�Rbm)$�{l�;_j�..����h�V��Xx�1c�ɠv��@b{̊92w3sf�77f�/�dLKˁ0J!�^e�5$�Ϫ3v(76h�٠v�ՠ^X���y$@̽�@9�95 �9h	V������0�)n�݄9�6��wa8�*�.���67<�%��Uم8��z,t\.�Q���� �M@9�ZU�1 8��*��+����O#rh��n��F���ء�s'��ﵹ$��~��9m��:�*���Dԋ@���sPG5 �9h��vJL�1!2�H�3A�ɒN���@��@v�ՠu�h�]M$��Rff�=��@jfY�����/vh��~m���O�v�\�gN鸔卣������|]V�a����W<� ��t����E���s�#5$��~w�u�hm�@/{f�v�N��id���@�嚀sPnj�r�&��us++wl �/wP�j ��GW�O b� ��F�ڠĵF�ABZ��)�Q��33=���;Šq�h��eI���0�RI���@�}�@��l�:�k�*��+����O$�h����sP䘀'I��tIt^�W�'ijsmu��v���q��ҡ��׳C�"y���8n<��78c;���o����& 	�j̒�t�.�/�d�
I�u[^���ă����/�Q�٠�u4\DXL�j8��5 �Ih	csP䘀�*޹��F,r94>��~�|������=�}��&/�x��4�5��SH�$+,CK�.��������������4Rb]A4�0c4i��e�<����,�s*��#H#&4�N=�]������6�f���Ǡ?��_�+csmpČፕ���)���M����y�SG�k�n�FK���y�ۍ��u �I�t��s$����zåxLM�0��- ��o�瘓�y�@k��4��"��gs^�؂��	$rh����*;�4����٠v��eF18�b�4��g�36h|݊ �fM�d�O{?|�\�>��8�H���WmzjL�h�ݟ�����\��&d�W�(

���;E��

��_�PU�AU������
���@cBT T 0T"�U�B(@T !B T"�EB#B#B�T"�T"�T"$!P�B
�P��AP��P��B�T"�B �P��!BP��P��T 0T"��BP��P�EB*T" @T �AP��P��B"�P��@T �0T *@T 
DT"
AP�P�BB ,EB����0��T +P��B
�T 1T"0��B1$B,B	P�,�0��B �P�
@T"��T"�P��T"0��BEBB0B	P�P�P�P�EB!P�P�@T �$�BDT$B,$EB0�T 1DX�01DXBBA`DT"�B"Ab�@X�)��W��

���(*�@PUj���AU�DW��_�@PU�AU�dW��(*�(*��1AY&SYd�>Y�pP��3'� a�_ Ӡ �t@  � @� ր����A�+��>�     U�    ()	 E��
�Q@  HH�EJ�( � �
L     �" $� (�)�})b�ū�M/m�\�_yꢁΞ�c���;�Zri�n�ez���({�ӗ_l�!�  �;뎞3�P;� (�E���_}��k��{9-�s���x=CҚ�h�zݛ;uEJ��;�  ;�TRT%(�.-H�{7���l�ۮ˵k���^�����D��׺�w{4|�:_s/�w�=և�� }�f��vx�Ֆ�`  �����3U{�}I@>|�j��3l}����y{���-����RU��3�����{e}��_^�U^ |%@�(�D�0 ��_qo�ԯ.� i�
P"Ԕ,�(=(Ģ�" ш R��l@�mJ)@�  �fPth�� �ePP΁������@R��ҍÔ��4ve a( �P D�@� NRB� T���)�!(PR��R�=�ﶛ羥@���ro��<m�7s�4�m�ޕ�z�Hn��;=�O.�x  mw��{mn{y�o�}H������5\{��w���U�3N��������#�'�����.�z�ww�� ��
���B}'�n�=���}^3�����=�r}ڕ�n��yzv{�}o���� �<=,[���N�  =���{�}��p�ܥ {�{r|�yy5�^���{oSσ�pu�m�۩�����]���:��   ����%J��h0CA�P��T��1 �=U*Q�G�L��ɓ@�i��1%I �@���%%)   "$!�)$@d<S�O������_����_�L�}�}�Ͼϵ��_�Y�TUt (*��
**��TTU�QQU���y�a�XH�`2����O����&�X�����@�����+�$`i�L�E==�2H�,B�P�"�p�)���E*�@��_@�F��"m<���� P�xM�����V%$�����>Bp+�uᆹ</:e5���}4�Z�֔���>YwOM:'���1�5��n��ZS��'�����fk�@v�h�!`H�4�����B��ʪ/!���`}*"�%]7|�Y�j]3,�l�s�p��i��`y$��2M�qP�ശp�߬�����K�'�_W�}��pī�U]]_���v��N�l�S���@�N><6�#�<�BŇ
�®��5�nGl��<���OIO��k�"��[���f�[.���G�L��<��k��ct�Zs^a��_������@������`��L���w�����\�k�}�ff��l����_��������	\ӳ��ath��HJJO���2�)��`Gg�~4O�O��hٮo�������}#����?{�&�=��w0}P>��q4Dڣ�i���8ǒ4t,
�Y�A����i��g�0��0��)�o�p#�	a^k�a�4��>���)R�|��A�"|��(�`B)����)M2@����:B>�=W�Lp=8�]$v{FN0��HR^<t��}O	]�p������l�|���]�h�n��:I��}36_mU��3����d5�8O~�����Rp��X��)=�i���eɢ4}��7��b|�$h@�53���i����X��J���^K�i�;��<}�{�����_n��5�0���!n���G'���ٳ����>2P��&5N��	��U*��o��+���r��f�g��L,��d(�y/2��Uկ^r���Y\Z��z�
��q�y��T�����&��i��)��$�7�K���7y�vC�����������X�ȕ�� �3�<I\ӽ5�s�G���,8��
a�p���:'&��)�jI���$���ޤ�c�7��[#���rIE�k^{�r��<=&��22�!�k�>Do���!�w�sp4deU�|�w��p.���8�2���&Ç�Î�r��[p�\4d��O��xC��_s�xJCLl0�	&V�k��)/�<����!w�HK�'(j>��m�9M��c���4n�
yN맚ߔ����XK������3Î��i.ȅ�|�xo�8�=)�߶sFh�,��R��k���4l�����d�H@k�M7ߌ��xMҞ\�ɚL2��)���0�w����y��JoN�56k��y&��L��h�+�dna$#�,R���6H@�2 Aum`�1I�A�L!1e�L�>š���$4rv�N5����rq6FF�� �ٳ�$3[�5�/��r�&h��n���IB!�n^� K,׍ۣ�rM$.g<ߨ'���W�>t��I|>�x{3������ύ������a���#!���$$#RB����ןRc�cLp	����$�`>@�<40u�!�`�Y������#�a&�+����A�F ���&�@�XHy�
9	-�g�6p��!T�R40>6z�q���ٜ6�BųJFͫ��wB�&�ɞx30َ�&�H��[tH�n�7�n������[�A296RP�P��Me7!C.���W��ZO�5�y�熼8j��D<�u��.{�ĕ�t�b�N����<||`���77��9��ߐ�˞f���0�nO9| S���~�\�$0���P�T�ǂ��Q�"P!C�h��s<>�av^_HU#IM{y7�5�x(����C��M$���␣��_8�c��E�'��P��H��:_ ��l�^>�IL4l�9��!\�������pѲO3������,�$
f��j3��(����NBG��p��j����rWP�u�q&щ�	�)�Ƅ5!�E<5*P�'��+�W��U�m����(�w��s���}<$7���@���<H];��a��<	
�,h��Mp7�2�L-��m�S���	�%�eIR$��||��Hn�ދ0�h �����!��}����� jPɱ�wʔ�����(��U]�>���Wmzk&��đ!`R:!�B�~����<�nh�<�$���a6&�yG�4!d�x�����$%�qm��Wfx��0�7�a�Hz���S�8���!��,(CІ!ɽH`h�f��l$�I7Y$�Zd�g���i�m����Ro��:������=!#R�B˨�������o��Ó�d�~`G:��3�ߟk��Vx�ͼ�Jx��ẅ�\4�M�y��y���{t�>XRh�y����WHI��N�4�_���s������<�R�����u0��>]h:�E*H��K�F�54� >���&�iU����(gj�����-��|�_�&����	�#�Y����^L��y���Y��K��c�@��9��l>�&�Y��$0%=��ILR0� �k��x�xŌ�^�a!>	=��FC=�&M�4�I"����Q���FO�D�0��bؓRC`�0�ą���V�f���
B���&�.��b��Jޟp���D�9�|�rzI53����4M�lI,�桱�CH]��!�=��(C�4��.j�4�4�My槷l% R��Q�-.d�8��Ϩ�O�3�;ڮR�TR)K�(�|#$o��7P����3m�9�%�ֹ�=.W��ڮ�v��o|]��/��Ϭ��?<dCE}M�'��:X�"�!6@!���E4�MF��!�	��	#��H0��8�<p���xl����N_>�4��>���㇞�'���047^@�@��x���(bA�~����I	O��G��2B���k�y�+$���Rϟ����g�I�e�RY%�,��zF\I���m~@ Hp3�֐ �0���P,���$�u�'��d=�a	����B�L�>��$��Ӎm1�P���C���d���4tF:�1���~<�O2|h���!���.�Ł@�D�������xBD�$d+$NB�H�ptd�a��CT�d,��&h��5>��{>4��$��=/�<���7���� CnɁ�Yk���BDԡ�	�<d$��'����yj��!� �%-�ϕZLȫD�.�dO$&,&�.���������U���}�p;��3O�}�S=��F�H@%i�5~@>����~ϏkZM�6 �jB�;�c#"E#�&CZ�9i���/�|�=�$u'�5{C��d
�i�a(�:<2��7�pq9"��[%���o�J?*��Gd�$Zl��	�&��Y�a��BaCz�!@���@"a��`M�<y}��� ���@Xq�RID���=%�����.sJ��#R���4|8�0��
jG��, ah�8C	 �觘�-C
�B
�
C��]�����)�'�R��!	�l)	,* ��()Sz5u����*�*���)�p��M!a��SI�]����
N����5GӁXv]��k�A�$@�>��&��0�$��_}�xi=��zCS��{̦�l�z�������G ��2lE�� D�$�K�������"U�O�c��$`���p�M����6&Ǉ�O><�y��n�[��
L� zH�.�̗V�L�*p�����T�� �g�
a�9�t��.���=���Y|y����G��S�Ov��<4h�8�{��9+��;ܗ��L�F~P��/���H�$BHf@�@����OC����x:;����,w��L�H	i�f�ӽo筽? �	�-	;"Km$���[[m�� �fݶ�[��i���m�a�)d��$i��[Kh��M�A�n����c� ;d�ֆ�v��]ue�cf��\���Z�h�Z�����[�Y�녹���;n��֗4Y.l�+��M��'k�m�m��ڻ�M�o�ݱ$�         ��kZ�   �                                H                                   � ��                   �    ~� � m       ��   8    �     �        ��}h    $    m      -� �     �               �   ��5��uު�m%�֜h�N���m� I�����#I���u�l�"S����H�V3rmٶ	   �:]s[%'@[@ Zkl�|��qn��m':�ݪk�9o�n�v�hͲze�:K����{[�mr�nZm�Z�$E�`�Y����m��f+`���:$m���d���6�.�6�I�!����� 	���Q�JM%ڻLJ�5������`a�ͪ���]v��]����k��́����2���i3tɵ�M�$sv�b�]��:2.v��X�8�̹��>[��խ�����/jֻl�0�u͋���` ��j�@e&ٺ6�ˇm�f��8���<f����u�mEX��lnԂa�� m����%�jV03�L�3	M�"��eb�V��*�݀    m    6�    �                        $    ���                 @ �   m�   Xg                                         �        �                                       �                                           ,7�e�`� p\�v�m��   @   $    m�[ ְ      6�      t�m�H$y�3�i;l��+n�cSb�vu��m�u]]m��Gb��`ڶ�kU�u�17D˻T�Nl�I���$Xm9�od#�m�k�l�v�5�ڦ d�뚍����L;i�r6�%�;^���$	8  I-d�n���5��V`��B���m5im כ=����l���`[v�*��4
����M4�e�۲�m��ճ�D�6�i�h��.�X���m���t�Y���`v��\ZY�M�5&��*j��B��SJY�G5��M����.�Mv]�b7m��ζ�p�����Y2�_m�1a�,n�IU�Mt�&H�ɳ�ScDl�DMI�r��8C�n3��+�[v����ԗ6]��ֺ���f��8�F�  #v��m� �          �>         m�  � �        [@      p[@ ���N�p�����ͦ�rr��gM� Ej�v`!|<�y���ͱu����U䭠:�..˓�&J 9"@-�sm�țΰ�@�vͰ�I4U�n�*moY1m �l�]0xK(����[R�!Sn�l�kn�h��4�Y���u�.M�WK�ֺ�Ʈ��٥ֶn���k3vK�XG@7 �k�&�iom�����2m�����T���iν����3n�l�Cm3]�4���]�X�3V�T� �9.�k����f�$���e���ݐV�.�Y���k�ia٭��II3�����t��\9�M&n�RΖ�6�@6�v�5�n5��˯--v6�Z��Xck�Rr�톷��`kM&�&�
�5���z�\��W$Ƌ�v�6&c�Ȩb�Z���$L.�Fme��n�k��M&t&�3kV�e�BEt�ln�7\m��ZOM#��ܷm%�B�J�]n��me��'`z��*L�1�L;.ų-]`Z�b�� ��l[�vٰt�In�l�2[:�l�(sn��u�ݲ��9��f�2"�[��f�YR*��Ue�b�hWm�h�"iYrIԝeЛ�ΓmkQ�\�d�Ʋ��u�v�4����m[9�L������l[*iA�ˋp;lv�f�-9��#k5RM�6i3ڭ� ?����9-r�j;2���m�qvXݸͻ��ޠ�N�d��OF�ۤHM�i:^��صӍ�m�2�6��H�\�54�����i�A���6�bp�i-��6Z$Y-�lY!��lql�O[Cm�j݅���J�Ip�ڐ6� 6����%�lH���-�۶P�۰�h�|8� � 6���Ŵ��y��  m�@k$�ձ'	��aq"/$4��\�H;��@���m�;�cv�d�����a�s��U�&Zl ,ڰH�V[@�km���V�h�u�ŵ�*�s\���Z.��z�H��:rF��]JL��[n��ʱ�;L���h��l8�[B�n+M�eL+�����Mש��ր)�l<�(浻j��[@�n�y�K4�z��۶���J)BM6d�:�6�۵�e���M�A��*j�,�i�n�	m� ��Í��Y.�rms��Y���-�H /]n��+5f�t��'j7d-[���Ŋ4.�YF�]�u�ʀ� Y���:�
�mL�u��ٻ6��Y&�M�V�&���� ���8�u�]��5�f�,]�`XI�Ӆ��o���m@h |>�w��In�u�޲m�;i�̰Z(n�6]����ۛg]r� q�Y$*ĳ4��6S��`��n�`F��fI�cm/K���]��-c�eC�����փ֮��"1f��j���[E���-kjڐ�ؽm֭��LĆ���t�T�N�Mjj�l�',^������n�l��ٲ�� k���[hm�l6�*M�Ukl�6�>﹵�j�m�1��u�� �i6�m���e��U���5�l 4��nS�Fچm(6tm�����;{f�M���K.msL��ٙSm�$-�[� �f�Mi�K���f��lؒ���M&Ü�&�$-��H��Xkd��K�.�M�A�k��� A1J9VZ�1[Sl�m�Z��`��9&L�ݶ�mIΗ�ݶ	 ��jmj˰Hۦö�v3k��B����� �6�I4��۴�U�ִ��4
bm�[%m�eY[U5��[P��W��4�6�b���]����t�kv n�7&�	ifskP\��Z�[gH�Z�[U;`6��8��Jګj]�l��޴�m6]�2��lm����:lZ�T%�W\�j�b:ٖ:i�ғm��U��bjki�m�8<��tE��ͭf�#Z�d�r�s��H� �-��Ͷ�Ζ�lA�V�ܤ-�vu��,�-��An['&v�"�^k�0m��� �]�%�n��m��R��t�5Ĕ�i0���u�p�eEUWm��uP�M/I.mk;Z� I��H$HM�6�ڳRK��Nf�vI*��X�`  ���1�]@�Xv�n7��kM�k�f�bL 4IV�*:Xkh +F¶*۰�� ����I�n�ͺ���/�����@-�l�.�[L�d�l�-d[v� 6��0�Sa5�6�:i����ɀ-�ݤ���&ն���۷�ٵ�"�3u���v� �C*�"e��`E8���I$�-:F� @  9Ͷ�a���g8�K�$�m�m�k�h p�$n�Lֶ��m�Ӡ  �[dNKD�v�F�K,�&�ۧm� ����� ����DV�����vݒm�Hl��s��m'N�C&ۭ����춶�:]6-�[8rkP����m�6�\%ՙLI�(Ql�l-�#vu� ڦ��l���ڈ4�}]�$�l���lڮ�֎�Z�T �b���@,�m�22iY�V��u� m������&��B����e��M�M���m��BKu��l 6Zڤ��lI�#���[��b��ɶ�$�6l����][�\a�3�$���] ��[w��t�Ki���m�Hl�\V��aq���O��n�I�^�W$�d�i4�i�jh�7Msn��6��6���e+��e�B� h�.�&ͤ�(�[4��A�kl�.����n����K@��芐٥4���K���nv��*��@�7�
P��1�cY�_(@�Ų�U��M���\��j�  6�}�}��e��MzYp�o����@]�_���CJ�t
�?��!�p`��"�#�*"��_� (�܁H5|F���!��>D�j�Z����(/ @� @d$b�OPڡ�<|UE8���AИ��* ��@�>�PO1d��'��v����C�) к�"��b�Q�l�+�#�T؁�QM>�!�	X)�: @��D� $��`��!	&#(IR#!�AO<T_�R�(�AO����!H �� �;t���c^(C���0 ��Wb!E�(�z
���@D�z0X��'�dd I$������!�B# �6xŊ�A>�M ||P�
�� HR�����<D�@H�*x���=O���EB*U��
)� �*�S�EbD 0$��m@�W�+�t�@��1J'����B�b�(�l�V�I.�N"��)8�>i�x	��{ وBz�W�R��dQdc*kD@�Y �(z+� S� S�Ҏ"���p�@��8�*TP�@M� �*��pTҁT��m0!P�D`-�W�� T"T}D&�xz�H,<L�J' ��] $@��@	�F*���3�X AH�U`���	 `0"1b��N �j&�^� DX��B��ChE��qB�J:�DbD6�(�QQU�G�(� E��) D�"X(��[��1�(�)�K-��"�
m�p�[�c���Z� [�am    � ��    ���   hm�I�m��  6��m�[Am�� �` -�o\��u���ծnufE�e�gLl�lX���itc-�R�ΰ���\֮%asK]��6��vօ�`@qh��uԺ�eZ�#�!3ir4�M��� �    �  	 �@[B@     kh�P ��      m�       Y�m�I�	 ���!m�f�[j�6��9�Jt/I%'��\�鳒/$'GmͶM���2�;\һlS5]�0)��3W\��#-��6$�^��S�r���  m� q � 6�m���5��u��-�4��(��Mą���l̶�̛'K�	�k�Hs�v��ėn��G1���Ҍa�6��"+���4I�����sw�$��F����9�&��͍+�n��.Я4-�M vm��U��qE�p$��$v:[]Բ3d��]']h����đ��}��$)zdלL����R�LT�Ȕ��5ũur��c�]�K]�jT��jf��u&�����˵�ЎK��9ذv�F���5�if�[��riu����V�sI�L��J��$�nκ��h�J�Ѯ���Je�M�Ds5f���ڲ�ve6G���Dt�f�vV(SM���V�r,q�F�T��,5�J�2Ԕ�2�n٣���t�uqs����7Zl$���Xm���K������Ei.ĥMy����M���ۀpZꀶ¶���YZ.͈[�-��*b��me��)�D�	��M���jؼ�E�8P���n�K�a(����P��6��ce�������Lr�4V�mun�YM��-�M�DԖK��\��	kh�F�@�Cl�]�-�[��
�]6e-q�.!:��/gN���F�Fp�W":�J�jf�+������=��w8+�A:�
`��OQCj�At�O�"/ C8�dB!	�CJp4����
;�6���;�n}f�L���f���tl��z�$�����4�mƭ�6[Z�����Rɶ�D��he�d�wS�vSv!L���XLʦl��\��в�a�˭f;v�l���ceԳ-�R�G-n�hfT�T\�IMp���k�c`ͳIL1��n�ں7�Gmzs4I	�3��cZ5Cd�2��т�c����f����1?;��UؼQ��$.[m�I�r̶�e��v���l]�ژ4֝a�$�Co�#���1�h��3�@;�w�{ݬ@y��GzṶ��E'#��Xו���ri`ori`}׺��"oiĤ�%EIGQX�� '=�ݒZv:��:Q&��DeI%n�����`ufk�7�+U������Xn��Q�P$hRA��1;K@w=�s� %�}��.Щ���c���*�r�t�0�M\��;lWJ�T��1�Y�l��.�Gb�� 'c�h�@N{�I�	�o%4���J���*+3&����(Cb�(uO��|����f䝾{�nI�^V�{��B'nqH����ɥ����g��K����ݞ,�$V�Ȇ�)��,��z�X�4��/fߋ��
^u)SE'#�	#@N�R���s� =rL@G6���1����b�+-���Σ4h�S+(�0�]qKa��m4��"l~Ȋ]��d6��r���� '=��$��u�fћM�$T�m�XܚX�& 'c�h��.�*e�u�V�HФ�����`o^V�Us��UN5�K3~L�S$~��]���c�ա9m�a�UU/d��7vx�7�4��U.����7��Z�p�W��f����@N{�I�	��U��W*���ԁƅ
j1JQ��A��M�����b,�M�6,l��4�.�h�8�s�E>ٳŁ���`o^V�3&�r�sj�ClR)J8X�& 'c�h��9�;ү]JT�I���H����`f��Y�r���U7���������I��ध�F�{���rEH	�`�w$���j� +�\H�b!h�S�U#ו�o���$T�swi9�䘀�����R���z���[a�tö�L���9�:�����Ѻq,���c/d�Bck
�#�6�B����7�+U���u��ϐ{6x�;���CV�6�q�G��yZ��]�$T���nL@IR��˹���]^�a�[h�*@N{�& 7�+U��؁o!�78�nJ�7�`�v���u-�EHt��V�b�H*Q��ś���s��=�k��/wiP���t2Ba����1;����V�y׫8����6��۶�n�Y+�ںXӍ2K7V�ԙK/Q
X�2��j����[@���ͩ���}��|l:��Մ��]3qZ^�5v��� J�[�t��[X�-y��p0�l��Q�D!K��B�@�0�j�4��VK�4�ۑw�jE�zdX6��5
��G(1XSZZ�f��m�����(n�b���k���$��ߓ�M�O=m�v�4��f�JKaaI��飍���0�sm�I\�B�i�	�kF'#�#�=�+�����XܚX�u��D6�ӂ���A(�+��J�$��m��@c��P�ZǠ���M�$T$ӕ`ori`b��`o^V���u`j�6��*���#B��ۓ�ԴI _\栀�sE5bTӑ�Фv��j�;����� �Ɉ	�����Mϲ��-2��#�ҡX�K�k��J��/;%��P��T�RR�JiF�*R�����,�M,Y��UU�c��=����q��*7%��ɥ��mQ]�\p(�%D�j��Шb�m)�COT8�j}u�3rN{��]�'�}���V.m+���AR�,�v�u-Uv\�P�����V��"��ӑH����`��������{���r*[I�JrQ���32hI&m̭?��@~��O@~|�qFܝ]{E�����m�J�	c,ٖ.ʚ���.�,�bjۭ%�.WK ^n�{�%�=2J��%�1WM�i
���HФ����U��ʫ�lJ����VfM,��5ՉSNGQ8���Ұ3^��TQʃ<V�������f��{��ݭ�Jikq)N�r���wZ��@9�Z�$�@N{as�6�8��n;3&�k�V��iXn��clBcM:��jJJH���L�*�i��j��v&��s5!�LܗLw��)��>z�U����V��=���7vx�=�s�u)�I��ȤV�IV��P��̒��n���b���@RJV��,̚X�uXkݥ`�fƓDtRs��L��2g��Ҁ͍נ?df'��fJ��ȉ#")2)��S��[�Kt�֐�:J�%$,1�@y�h�5��|�pnZ�Z 9[Uoi��b�Ƹ�1�A۫4�����]i�mI��f-����Z q�@s{���H�-mȊT�:m�V��/�+��$f��`o��Xcݥ`ndT-�qǺU�nf��� �-�U�3e���*�W(m
E �,=\�s�ѯ9�@}����//&�Y�2{̭(k\��Jn�Rr:r'��=�V��4�s�y�@��I�F�éQ�n^� ��n e]�@�uqh�bī�3��]u��i;nm�t��LZ�ͧU�sm�l ��w�l�ˬb�ю��^��$$��GZ��'Cj���M��l��F�n3��m̦,F�`�Y^;��6���6�e�݊0��m����k�f���	pmm4)���J0SL:ѷ��o��CN��ly�;s$�h�S6��5b��t�t��|�����w�Zx$&���Ʒ5!�Й�X�-.�Y\d�����Ԁ(��0�Y�V��ڿ {����o`�q�y%Z ͣv4�":)�ErX�M/�*�������?z��f�˾r�#t�֐�:J�QHXܚXu�ҳ��F�},͞,��f�QQ)��),5�?�;��76h������#B֣E*R�6�+ �͖�\������,��iXݥ��%C�_$q��ms�B1�,��Z�#�c�b�Z��`�*T)�4�B��ܖ{�Kǰ@{�J�_}���jҝ����)�����ɥ�UmQ�Ts�$a �D"�)�W�Wۃ��U�$�s� #��L���B�������v��f���ɥ���K;���C���@�$�`9��@8�vIV��,�4�":)�ErX�M,ܚXu�Ұ��`]UW�M��i�H�EU]�u�P+��K�"ٜ�ty,�!7h��4%��J�!Tt�	����M,��E`����ri`}�36���M9mH�`}ך+�$���36x�3^j�W8���R#B�Q�RR�7 �}���y��n|x�q})B�F��������F�������# �`D!I<y%���>:����x����rs\<�$� �>������ˠ�Le�$db�C��P0�z�	�&p�a�HD�H�n�%~�SI�%+@��Q���x���p6�cP������6�r¡�40��֘,aP�"�"���!q=� �hš�,Z�C� yu���R�h��������q�6�2"D�,,f��&�$��ܗ���6q�Tt�����o(K�9#�'�0LGXT'9����0�L5M�*�*5M�M�H�ц��u���M.�CU���(�]�z(x��SBUU�E`@؆�\@N��z�E�M�^�1�hLP��8|� ������8��G�g���rNy��_��������T/܃N8�)J��a��q�o�(��z5'�1k�bd��sf��tg�Ux-��ФR"'|���ʤ������z��͞,��xlksJv2��K1��t�3��λ�j�d�׮��Rj���0�~I���i��-z�F�����d�~s�}��zs�ȇ�虔L��O0��<�DooMy����lf���h��L�(�����i:DtT�ErX���=\K|�^�d���h�y��� �ޚ]aˡ�u0��L��%s3s3DѼ��oS��2w�krl�xV���
�-P�(<�*1 �E�B�z(z��f~�����d��'��MSNGQH���¿ܤ����36x�ߩ�-�wk�m�*�.��p{b�դ�e[i{V�řh�f�lİ�&�R��)4�F4H��Jt۔�ަ���~�o���QѼ�I2�������nˡ��i��)Q�,��{����y�������gr�l��(�D˼�C�IAɗ4vV�������\�7���/6x��˒Q�N��J�C�3*f^%�|�Q@s%�=�y��y�ɹ7��.D�*eL��̨���fnI�2e�����w��&o$����ܓ�o�V�E�F*B�(ޗ���ߚ۵��ڻ ��[)s��d�nZ���x��e��A�l��&�u��K>�|�[l �d`��s��ս�lj�V��2�Ѣf�76��Iv�a`h�1e��p5.6���$�E4�vlWB��X���ݍB�NΚ�@���tV�#�\�X��4i�����m0�#(�&í�l�^chZk���D�r�k"�7e-�;Kc�g��}�I����	�[i�Ζjeb�+��Ki�n�0jk�m��f�Z��j�@03��1U��ra
dR�3�̞���͌נ=U�y�y�	{|�U�kZB�:P&�EMQ���z�$�k���K�oE���jL�ϭ��B�D��bb��^�׼�(ԓ;��lP�:Pk&|پV��H��h�%D��R�Ź����1�@;�@F���}�\�9
R�rXܚX��U�����|; �͖��Vn߁����u5yMV�6:��P���n�˳��v� lҹe���r*��&J�D�`�:����w����t� ��L���,MI*H�VWsGy��Wq��)B@�������?f�{����\��tA��;��*@&���~��`��7^j�:��;V�v4�":)�D�q�~�Us�7������>���gȋȠ1��,�B�:P#q�`n��`~�������~v�͖u�ؔ
N��8IN��Yt�,M�q��8���U��a43���cX�f��FwEED�䍥��5f�v��v�͞������W�D4H��(�w�"���ȮL���ޚ�7�������Ky�q�R���ş}��{�{�܉��
@���+��@� j��w���~�ܒw��[�s��0	DB&]�bb"b����̉��1�WE ^^M33tl�tP���
St!5$�"qX[����q{7��3^�Xך��)m��	��u&�m��役��V�\$��Κ�`gB\m�l_���ӡ�I�Bi� {7���<�`o^j�*��[����=��t��Q-/2�3@gј��.d���z�{����k�&nd���ΰ���:��F:�B������՛���I���=��Vp)��TPI9#iE"��/=�"�6�f�ϣ1�-2Is	&hd�����7��������V���P%f��9�@~��������܆ ;��B؍4
���@ʃc��h��*̩�h��G��xKsI��҇�/�sp��a)''�{=<Xך�Y�?W�f�X���	��"�$,��W���S&�5�t��w"�ϲp�ffK�A}�ХD!Ǉ��3/�>�@~|��9�2�;:x�7#y���� |P�%'M	�a�]~�;����μǠ�e�ӽ�P�t��	�(��S.;{�K�[�|��}��-�v �b>�}>殌.�L.�k6����^���$n�H��9�T�d���r����)i��;g���m hZ�nF����K��ٚ]F��+�����s�U���-�c�)k&��Y`X�+��s��Q���5pQ��f����CU���FT���mYb�î���0�kvշ�3�Gg6t۲Ռ�M�c1v��Qyi���tΰ�5�9c�:m&m9�O�I�w�䏯^:���[a�_���m���R���2���K]+�UlZ�\�xfIt&7�H�_'�)���-�i�F����E���?�7$�&C2_Hvt�@g��
^Gw��r�����Ek2w>}͊ogJ��ǭL�͵�CĦ�TJm� ��o���٥�̓rd����>�4���wN���B��!Jq��K��5���InM���n�ZK�UM�{|��$���ui�!:#�����K;3W�$���W*��xs�$�����$���ZI%�,�؆�f��f�Ju�����t���[va�ήa���nx���>N�9�Fm)L+2~~ S߼9i$�{���$���{������/�I/{�$خ��:hM89i$�{���>E�%�`(.)�ܧm��KI%����$�����6�^{ѧA�Q�*����$g��i$��{��/�U��Z���L������9�m���֐��J�u����UM�^�}�I}��I%�����/r�+�{��Ig�c~{�#@ʗDSנ
~��W���g�ϽI%����Igfj��]�JS���5whf)i���Ԍd�vY2�5�d�͝-J	h�j����y��� �K��|�K�����$��b��Yٚ�ʯ�+����>������ >�p��`�gz� ~{}���t����y��� >����{���z�;�Y$T��}t��`kV�9$V�K���}�n�ZU�r��RH? �D<�s���r�oߵ�Wv�}{���ތ��b�7נ<��O�^�ɪ�{��ww|��ߝ��윗�w�nd�;��翟�o�@~�hmO&�f�b��Mkv�y�{�s������P��߿��$�����}�I%����K�sjE���h��@v��B�p��BX�6mr`��Mr`�+5�%&MMRR^��� k$����r�GȪGbI-�?Ei$��z}�I%����K繯�I*鵭!ThU*2�̽;���u���ܙ���ɦe���ַm������[m��}����`�0H�T=��7��Q�h�t\�^��߷Zݶ�g����蟘�"��w���Z�n���ϧ�@粷�f@�M�-u�oT$�DMk�����-�����wm��5�ל����$$Z�X@���%.�?��W~k���Zݶ���� ?��\�ms�z ������~H	�y���m����5��m�{���[m�����P�lT�p���L�*�i��L���l陠մ�Ir�Kz��#tkxp�`kV�2(~ �?>�� �u���=�����!ﺶ��Z�n��������
�L�� S�߻�>t��!��fi�w�������:'��ww�����~�A ���{�d�va3 �4&���Z�����%�sEi$��5}�I7G-$��Q�#t��*��T�k9�oD�C_~�?K�m�w]�y�m�߾����!�,R��~���r�I��O��)�Zx ~~���^����.od%5��n����~����D�.�����`�J��݇��{�BW?�~����°�>�6M'�������ap3C���5�@�С��p�Ɨd�'ԡH�����	�$��޴w�2�!�s��sA��E�Φ</8�p�@�G�H3˚e֪D�of�K�����N��(0� �� $�Q�� �aA1o�;!�@�a�	���Ɣ���"�� F��
6B<6����I�k�����@�1$��ᙘD��͈i;'�$#�_��`D�|&��;�s|O(a|�y����&a|t]�,�CӉ	$��Q�f�O��hF: @-)�`�d++
h�R�$���Ҧ��O7�	�b�6>!�߾��/�`Jy#)�
�,�\1��y�pp<���h\׍��bCZ0&���P��z!LS.�y<�98�si\a���e0M6�QpwT�VX��v�+�JJ���hAc[����v��ma�8#��:kl�  [u�-�     ��8      � �>  -�mm �h  -��m�@[xH m� ��Zs�^2֙۶�GA���f�j��yMf�q,��l�70%��D�K����Y-a�3^�d�I�n�7,9����1ȑ��f3��l�k�Yp$@6�    8h  ���� ��  Z�@�`m                q"�� ��n ����"X�����#��s5m�b�m��&���wE��mR��irj�$��.�v4qL��9���&�-P`W0ՙ5(\�FF�T�p �i$�� �n6�ۈ]4��3-&�Z�©�1	6��ˉ%�!m3p۵k��e�(P�Z�:Ԁ��	��	]�v��v����F:#C�d��+bfa����ͬ�8)r��K���K���EB�eR�.����)6Ō�t�m�\Y`�s�i�ڄ�M�,�����ɥ�ڴ�m�s�m5S]lٕ\P�ĭ�ٯ�B�Z�٭���0��[�@pmB�� ���b% [B��l�u��8�y�d0%]`X]jM6��u��^e�\�݋����E��[�bV6�4�S.���4��M�m�ճ�{�����n�kq�L�.�5�L�\Q%�4\ٶ,���,Xh�xR+
�b�[��!����N���*�&�t�8�h�e3]����Gkt����Sh�խ��b^V�d�:k6�u�E!%��m�Th���Z���M3U�P�uvM).J�Ef�ZckqZ�e��E���l3q6�K���t���i0-�B�	�e�66�]�k�JWWk4Mz溘�XL۩�,s�	���:�\�]�K���H�Yx��f&K�iГ����$��"^��6��b�Qp-ƥЛ-��+6U,3W����rh@�Td�!�) h��<��  O�D<}E6�mJ�@8��T�
���'I��߻{�:�i�����5� 6ٶ�z�}��]dΦ��Ζ���j#�8��h.�6�WͶm� [@Yv��^wM�l���W�� �gET���,vk�څ��[�m�XJ��n�۶���th�1t-�ٍ���[�q������l1�c\+
]f�qh���jDH�ebB��DcHSb뒻m�fD�cf�Ɖ��e2��Z��;����H���. sF������oXC]5�k�+۫4�/�J�u���?��%�Xylo��H��R�|�O��|I%�����%�sE�~��-�����$o��f@�M�-π�������뻗��G�ߟ}�����'���;��y�M;��̴��A�r�G�$�u����L����+�
�H/~�9i$������%ݞ���WP֭�dZx�>��}�����-�^��3[����ﳜ�� �C�}���� }���q��6�aX��נ
~��t��_�������1$��i$��5}�I/����ZaI,ѵ��@v2Ć�]���6��<�l���V2�B���>N��񺎘�0Кps�]{�?�I.�+I%ܙ��s�HY�9i$�u��eG)T|��kY�[o�f��]�<|9XD�KN'�8��y�kL`���"�ѷzM�$!���Ģq�����?����;���������x��ww���y��7/�{�<)>_�����������z?~ww3&��s����ߝ��x< ={�7�ܩ�*].�����XTs����I%�~|�][4v��_�A&���������3 �K��93�������٣��]}�|�B��夃���=�	uƚ��\-����s��eC^Y]��h�P���Z�:�p;�:}�'���=sr��!Jq�$�����$�_w_�$����>fe��ɒ��w��z?~ww�/T*xCZ�)��x ~o�~��_{��ܩO߿'-$������Iul��I,ݷŮ�7I&�� �|�B��夒������18�W�� pX&�N u�W� �"@�		U�r�����}?�i$�=��|�Y�'�j]2�(DDK�ӻ�&�/$�*����~�m���K�m�g�}�����X�z�ߦ@�����5��;�ʾ� ~��um���A";�;���/�߮ki$�ۻ>�$���= M2I���E]�u�P+��u
�g4]K�Ifհ��Зd0S��B�:H� �R
�IfL���$-�Ni����fO���̐�d�N�����|�lo��R%4T�c'�@��ٟ>�.L��f]���k�GOCӻ�������O�[�gUC�ҿF`	v�g$��Ig�ߧ�$�^�j���Sovo��$�>|�/��~� {�s��r�נ>� "�o����.�����ל��~��n���Ƒ��-ZFB2$�Ō!� X�0�F��� ،4 |	���T��Tsޙ����$��?����H9$�]�m��{��-���?���M����I�$��������٭ZI,ܫ�@8٬m�J#���f�e���s�[��˷8��Ҭ�:Y�ƺ�Rk��ћ@0�P��� n��I}��W�$�u������Q]�%�O�O^�>|ɾ�QҊb�d_ Y��~��Ʉ)�|��ON��;��󻻾f���l�^�P=�/͏�X�#����I-��]+I%�3W�$�[����_o�~��@��`�b܊��?���'�"S���������������m���s�ޡ�@����vڷB���(�Q)�:i���$��-'wԹL30�!&��Wn���Ԟ����~���m#�Z�c�I�$LG�[�D��w{���ѩZ��0ź� ʆ�.ܹ�Kn:)���-Sz\�*i$Š�l�kp�vm� [A���Z�Z�4�,v��1���:U5t�� Υu�h]�fk+u%����\fcm�]�Յ��5t�,[.M��01���K3�֨�j6ru2�o$��{7M:s�l�.��Y{s��*pisUF���:��)�hf�J�vˑ�#u�p�m��mְ�svڒˋrKխ�Kڥ��-�F!6����5���)6�Q�]��ȿ���p�-�ϳ�v�}�^�
�/� �"���e��� ��������[�g�@���!�����['Yb�������K���KI%���}�Iwi뱲AչL� ~�~�^�߿b�N��xL&0�Xɪ��U*}ޥ@~�'�2aM]j�R�ru?F(��#;����@~��T�rM=���S�(�"hhM�����u`yȩ&Ih����+%݅�����L�Tv&��շQ܉�6.�.5��ju��4�Ά�I��k�w&�V��6���@fcβd�8n�Ҡm[� Д����׺��Uos�*��V��Q={���]nI��}�rN^e*�$˓$��Ptrx�%�S��^%�;���̥G$��4E��t~����4��R$�lm�I`n��P]�>fE&\�(��:h�N��;���Ȟ^"eP]�3&K�e�����4fe*�ֲ��%�!��o)�ۆ�^�j	�w�鳮XH��{]2ݲhe��5��ڭjܦvo��g�Ƞ׋&��̥����@f��@^t�?B�'D��yx�(��ɯ&Is$���Tn�fN�˨� y��M	�RX��Vs&�.W���2Tɒ�2�L��jt��[4�9q��L��a��T�&䒌������ ~�Y4�&}��ʀ5�f���C��H���������(����߿]Xך�����@�t7H��Jv��VՁ�lsi-�Y�61��� k�Y�o����[�M��%(*�à���X�����@I6���+n�v��0x��3@ffR�fe̒�/cy��(��ɮf\�y�L�O{����#�G�(�����+wf��el�7wn��n�$`�9�����I3�3Gw~�/ut����)/�8\d$$B$	2B�c��H�$�$�$���2^3�fW���{���2���n�o3D��L@I"������,6��l�jGQ��$oc�yongG<���	*4ٻB��*��C[6��[��Id���}zn���..Ǝ�����J���^E����I7!$��ɾ�ž���7�<�_�*9J�*1�V˷�^L�������-�32�k&e��'O��ޓ������+qA�q\�����??ֲ(�3$��wiP=��v
�O�䧑��IA̼��&M9�����@~�"�[�fL��@�ww�(C��1.�����EH_9�	&���SGl�a�!����_g��u�����,5�̠�m]�����ҙ׭��I�6�P�Gh������;[-�u�K&� ��m hZ��n�U̍��Yfa[e�&eSF˪1��X9K�6��u$�m5�����ۮcv���s�iZG��]�kl٭A�Ҧ�61[�6�֮Y��6Ѕs��f	�l�^�X��\fF�ܦ��"�å��j��\�Qu,e���Is.�h�s��߽'��֞MlHѳ@F]T2��f��+�
�Rf<5�ҰIsf�m����Y$�/Kz��&����G��nJ�����`n����SH�Τ�a��Wx�2�1@fd�_̓77�d�&C0&i�yz({ޥ@~�"�̼���d�&�o����u)�*�EJ&�`j���vvEH_9������M0���o.�!�LPy���xL�&N�޵@c�z(��(<̒�^Bfa� �o/E�{��K�����
��*��w5�͂�Φ :H��ݽ��p�5��O6�x��*��=Yce3�A*dU�m����̒aL����a�xrC�je�F�WVfn0?����D��L@t�R��b��T5�M�"R���,�r���*F��B�KQ!2&a�ơYHm�&F(E| �D�2Z�nI	�!2OE��@k�tPy8W&dܙ�@ha�(����w����1@gwR�??בG�&L��fΔ�x�<����1��j.v`�,������Y8�fd�s��@n��@~�dPs�K=�}Vm{��4�$��"#�.�p�93y$3$�d+�����Ԩ�s]�f��6�6�N�Cr7)(�YiaI��E������n�Y��x����!R�B��R&�`|�������X/�#RK�L�>������u$1.�r�2�ܓϾ�f�'ሌB4Ao��@n��@~�dP���>@
9ITM9V��U���K%w�]�Z`�����z��k��	|�O�솉y�5q� Ą`�5����r��H���<)�MVnM5��^cm�g�Q��C�`Fv|9Æ<1�M�����R]�a(F�&a�.���ej����K��#Į��X$��1H�Ӝ�b�6|!���ny��@�z]>O:�w�/ړ�����F\J*F��p<��Ѱ:_0<i�6h5&�� ۰�1�{��7b4pq\p�H��,`���
h�Fh���.�4��o+
B��Ɓ�����A��,��S���ָGSxVb��#[����D���j���bl�$�=EO�v�iF >��qCb��=�_P0�!��� ���!�>4> ���
UT*�PS��V�����7!��J�1�X,rHw%LK��̽�$��6��1���fR��oɢ�������Rn�F�`b�V��������E�̙�u��k5�eS[��% �3g�W
�k��fi#�Q�Ѹ4sn>t�׻�^�Z�/���W ku�%L|wu*�E��y8y�3.Ixd�HfW!ϼ���uh!�bb%<������- �� ��*_���/K$���>��]q���(d�������u-�"��9h&��y1	�Ï.�1%��&hܭ\�}����9�{�ܜOP�m�
���L4�!�����A��B0��7.�D�l���\˸&(�lVD `U��Z�ܛ�w�����EM1&'QX��ՁꪮIy�ff�~�=����@_�k��M�����n��Vk�2��j�Yj$�P�2͚�˦�D�:���.����������s�_[��G)"*�7+ ����X��,���`w��V����DD����d�Z�a$2DA�����T�p�3����I�DJPU��޼�V�fR���e䆙����7}>(����rD&4'*+�ݺ�>��,�'
e�J3+W=����h�&&"U鹻Ht� ;��ݎ��;�T��c��cT5,7�J`A���#F(�`[QjI}�����8��A�UU��*��R���n�Y+��o���a�2[wV���K1%�2������V� m���I��.���-��t�!�F�tQ�BT����B�3k-,,5),��e-�뎜M�Nٓ�I��v�4i�yz�j�[6�B�`��ʺSVZ���ź2�0�cl���Z]�v�h�12bۮ�b],]�.08�¤�b���n̳!u@͊��4��g���z�v���چ�`4�����^	�eZ�]{L�䩙v��u���0����<�z�i�I��D6��=����;ו���wn��s���;��,g��^�ҤТ�jbJ��=y���_wR�/:x�.�p�3&KɓxCL��Q� �"e�<x^V���Ht� {_:��;��ְ*9ITr�=��ʠ�qE��ʀ�����ZȠ?e�* ��aZ�4�Q�rU��ɥ���_���I!�\殏��ޥ@~���q`f���sV�V�[�ipbZ�q�a`f:��@��IԞMn��#�k�ٿ�����������^R�&�I0��͞,څ�ȥ$�PhnTvۛuj��RBS�`V��E���$H�!>A���ٿ��T^����Ek&f�K̙$��=�JxH�L��y���@f��PܚY�\�K�6���}u`w7]�jH[�f�Z�5���@?�2 F ī��>��P��H��@_�0���!	�K�K�Ĕ���E�dܼ́2F{�j���R�/�(�b��e4��"DI�Z��9z�L:�!�h��KY�D�tՌ�7[�k@�be���K�4w��YyJ����*���R�_@[殊 ���k�9ITr���u`gri@~�dP��o&�����$�rT��<<ʠ76x�??ֲ(d��̄� ��#B �߻�rO���V��V�)MR��Q�X~��כ_�ߧ�Hs���� >�ܲ�[$�������X�w&�|��˹Z�̥��%Ct�JBj�lB\6�u���yev5�%�*��W&6��RSRA�Rq�ȓ�#rU��^j�3�4�??ֲ5��f��z���A28���ݳ/v�����S�*@{���W�ޘg~�!	�H�y�(������qRݎZ�� :=�ɤ0LK�x��OA����*r7�rO|�_M�4	U-��`(q���>�w$�yg���Hk4[5I""UE����B���|�o'�>�۫�ȁ�i�H�5I�*H��ĺ�R��[��U��]f�),ڡl�4%3L�5�4�Q��n+:�U����VۛkS70�����>��3Cʘ�3m�U�=T�}�Z�9k��I>Ο�*���O�Ń�VB�2�B��H��c���{(@7�����"N���V�Wꢟ���X���hG������1e�w�f�ː�/@_�x��ܘk������Vu�땙Odr�!QR�Iź� ʻ^�l�N��z��l�u͜o�e�'�]zD�Atٴ�m�m��������s�f1ڢܚ����Fܚ�j�-�v��m1�-�9���l�3dvm��p��T&ͻu�9#]/cٴ해�����X�l�k��h;;e��p�ʍ�e�Xp��y������ɣ�Jj�׳�*5�F�\�Ζ�5���%+<��۝��6�%j�᳞�;Tا����[��2�v�yX�fEĲ��m��tRuTIH��g��>�۫f�&^Be��o=���:H"`��Dy��B��Hm�@>�-�6P���Bf��6!ߐ)�N互"%P���� c����(@z8� O�@�rHw%LLû���I�.fd�r������P��&d��flP��jFƥF*��`}�6��+��o���ջ�`g^j����aI��#S��ݶ���+l�kݡڥ�ĬD��P�[F��\7�)��)F�%%�9E����X�5�ܚz���}��,ݎ�~��f�ִnI��߳x}(*#U�����s����}�|]�}��W���;��H!0QȂH���z�Fbz5$�2Izg=ޥ@s�y����E'PED����^�+�^R�-��(9�'˜נ3pO�'�&��e鷛Z��qR�s��@n�K:����4�i�@�u-�[�n��hl\�*��[f"c1�'O�d-�����$EPm��^��`g^j�I+P�*@�P*Y�]�[�{c��E��2\�@_w)�/��P�z�]�*FƥF*��`n�K�s�~ٹ��y��J0
F�:N�$���L��r_O?}�@f�s�z��YI"9IA&��,�6��ř��μ�a�\�]��R�������<RDD���E��ɻk�� ��`nl����m�m%P���m�7:i��-ӳj�htكn�1�52L
�\MM�Ƥ�(�A$v��V�wi�y8j\�d/�5�z(ޘg~�!	򴲶��m zIZ��EHm�@K�ǮM�!�Q���zR<J ��^%M��J���Ǡ2�1���ɠ�e��=�c�#����$���g^�;�y�t{�@��M�M�&C&I�/\A��_xnI>}>���L�h�j�Ľ��@y���a�I�;����{�V��U����"P8��$$��k�B1`G<��A�R,ś��i��Mb�h�k^E3wM���7t@n��'8��U��ɥ�w�Y��i�J	ʎ�ϯ)Ws!! ID���n��̭vw*:)�������V��U�s�̆E���;;�P^dPƤ�)#���W*��oŁ՛[}�J��I4\��P�0���'Ȕ���}ܭ��*�\�{�W�ug���>��}7$���	�>�>t��O��-|��P�ٲ��r m�G�܏�j��@�<q��ޏ���>d���I8}���@���x��OD|��=#���4���GBx�v�9�A�������J�����@>����<����sq&�E�'��Xm��>L�<16<A��OF�7HM���0�$�7��;8:�6BMD�n���%������
�R�1�`p�H�w~I�;���z}xA�̢��e��j�`�u���	U���m�[m띶�  ���     h:      '@   -�mm �M� pm�@8 ��� � mg$��26�.4]�$fkyة!t35�Ceث2LZ`*Ken�p�θ��RYZ���e����p�F�M�n���1k��um�[7rS���H�     �  8ж�      l$ ]6 �         �      ��E�(� ,з [Vз%��I+�㝈�N�ɝΔ�%D�HI����3Uvm�.���۔�\�2�W]M+@.��;S`��7-��--w�᷂��Uf��]�  -��8� J�i �33-&�Z9s�V��m�����Y����&Z7]Dҋv۩fuY��tr�S��m%�7�c�n�%�Z�1������l+�%x41&t%�-�\��� q.ঽu���#v����%�4��%D�n�4LuvgZ�BrF�k��6��t���٭��۲۰�%n؎Rۘ�mpś*�h	C��˰-��XfR��u��\3S[Kz▻2�WUf�5M��ڄ�Q���C[�6�KT�T��PhYMI�x���41u��E.��F٭٥�s��mօ����j�r�ݫ�!hff��;`��ƭ��6m/-6ى`�K�[��&[�.T�-ɵ�CA@�F:F,�tꐫ�i�!����L�ʂ���^t�hU)*mI�Э�56�4��n �퉃�bX�\ݳ*Y����5LZ!�L��$�νd�Ov�W��b�@[Il5.+3[5���d�u��"m!�ZLL�u3�p̃J]����l�2ؕ$�c��Az�sgg1��ڤ�$mnD٣�^�z4��&BP�mUm�d�	1�]s�[�\�f˶@m���nM�4[-��-�+	ft/M�i�.�2An�Y�K�Bj�Y�[& ,F� |�J+�#����S@(|!�
%##�Ch���|Q �����6 x��1O�C�  >�3	L��\�N����@l�w[6�N	�-eS�����"���R�zβl��[��k�m�6� -����61�c�SQj�)i��e1�D]��2��Iv�%�&�0�l:�mQXMGk3��5�eG���]jV]-1�%����3��ыK˰�i֭���B:R�!�5���e"��Z��Kei���ͦ��,\����2dIF7B��՝$�M$�򋶴�0�:,U�e��E�hR�����n�fԡ*�SM��`v��-��i�q�3�m���J���^E�yK��7�����/��i~���$EQ��X.�s6����ZȠ3��U�L�{�d&S!���O�S����v����V˹Z���Ձ��k��V���H��G*��������o/E���P��Ƞ2�)Pu65M"H%��G`own����n*@�SP�LU�[u�١G0s��T0kAe`��394��xk�c���D����%�׌�����\�	��?-���@F��u5:EHrb0jA	���r;s&��+y�U}Ó����EaBB%��``B���3��i �*�@t��P|�fQ�!3	��w�]4{����������"QI�&�`w+e��fR��d�$�-�z(ݞ(��|����	9#�%��ݺ�>]�v�M,��l���[AQ�J%Q4�??ב@k.I�������h�6����ڑ@qr2�5 ��d���*��<��Xf 	S.V��v�m����$�^ciF		$Q��`nd��ܤr���ͯ;�|r�K������'�2%�b{�����N2q��Z��LJ�
dֵ���Kı<�~;�NC��DȖ'�~��Kı=ϻ�6��bX�'~�}�ND�,K����)��kR�Kff�fӑ,K����"X�%��{�siȖ:A����S����m
hV�&�0�)�9��*Xp 7���~���~�}�ND�,K�~��6��bX�'��ogt̙�l�[�Ѵ�K��A dOu�fӑ,K��{��iȖ%�by��w6��bX��̉��߼6��bX�'���925 ��H�9�9H�#��V�ߋ�r%�bX�g�ͧ"X�%��{�ND�,K����ӑ,K��W;���]�.�ƕ)�,@�����qA���7f�,Y��R����
VXh�ۮf�Ȗ%�b{�t��ND�,K���6��bX�'���́�E�șı;����r%�bX�~���^�5�[��f�fӑ,K����!���,Os��ͧ"X�%�����iȖ%�by��w6���P��ꦢY���_���9��v3<���/B�"}����ND�,K��ND�,K��㹴�Kı=�{�iȖ%�^���{��͆˕vw�=^��Y߈bdN����"X�%��}��m9ı,O{���r%�`tG�x<r'�}߳iȖ%�bS��N�Fc�Z�0�f��"X�%��{���r%�bX�����Kı<�~�m9ı,O��xm9ı,O���K�3�`��5�ѕMnT6!��c6q�%p�����sr��C��ڹ����,�:�z��N&��Զfh�m=�bX�'���m9ı,O3߻�ND�,K��ND�,K��㹴�Kı>��xC;�d�[e2�֍�"X�%��{�si�
���j%������"X�%��w���ND�,K���6��bX������ޮ�ZRasn]�OW�z���ND�,K��㹴�Kı=�{�iȖ%�by����r%�bX�{ۼouf�\5I�ZѴ�K���`�����6��bX�'����iȖ%�by����r%�bX�����OW�z�z~��m>kQ�qC9��m9ı,N����r%�bX�g�w6��bX�'~�xm9ı,O3߻�ND�,Kz��F5k:��Ν/Y'���;CCBe+a����S:�k4�u6ͫj��وZ����9��JRɶ�D��h [@�@ֲ����]�+�n-%e	�fv�7e@.`+5�ZScj���MM�I��7r�V��iIs�X�չ�A3��c���`M2�X�Ͷ��i�����W9X�s5�5	NKS-�Q�R�&��[h�j�aCf�U����X��r�bgM�t�Z�j��!�\E���O�(� ��T�/��|52K���{$�*F�[m�E^�RX�6Q��bk�.�1���q�kiCv�V�1�맺�%�bw�߹��Kı;�{�iȖ%�by���� �"dK�����<���/B�/C��>ZS��eʎ�|ND�,K�w�6������W"dK����iȖ%�b~����ND�,K�~�6��bX�%=>;d�f:5�35�4m9ı,O3߻�ND�,K߻�ͧ"X�b؞{�t��H��v�3 L�����܈��ʁ$?@�U�?D����m9ı,O~��m9ı,O~�xm9İ?�+�ފe�d�'8˻Z�
:QK�)��jm9ı,O=���r%�bX�`A~���O"X�%��}�ٴ�Kı=����r%�bX����fj���Qk�e�β�iq4Q�E�.Κ��b�Q�0m4q�Z�,�����Kı=����Kı<�~�m9ı,O~��6��bX�'���m9^��^���y���)j��ŉbX�g�w6���� �T���P�~�H��"{�����m9ı,O���ͧ"X�%�����#н���i�Xz�3��]�OU,K����iȖ%�by����r%�~ B	!�2'����ӑ,K��>���r%�bX���2޲kZ���W.�6��bX�'���ͧ"X�%�����"X�%��{�siȖ%�b{��iȖ%�b^�>���.�3Z��L�fӑ,K�����ӑ,K�d}����O"X�%�����6��bX�'���ͧ"X�%���$�����m6��ah��mU���5)V�&�Ɓ��dv���[m�R�y5�1�,�L\,��Y&f�\��{ı,O����iȖ%�b{��iȖ%�by����O"dK��~��Kı;��\����f�����3Zͧ"X�%��{�ͧ!�b��,R1��MD�>���ͧ"X�%������"X�%��{�siȖ%�by�n��L��l�K�Ѵ�Kı<�~�m9ı,O��xm9�K� i{��p2��)hJA�	(�j��1���z�A�@�`G蝉��s���Kı?w���#н���ϓOWj����ۗy��K��H����iȖ%�b{�w�m9ı,O{���r%�`~dK�ފe�d�'8����\�<)���kiȖ%�by����r%�bX�� ��0O�~���%�bX�����ND�,K��{��"X�%��'�T�2���+-kn��$����I)��f4�a��%�V2��n��]m`ƙ�&k5��m9ı,O{���r%�bX�g�w6��bX�%���[��DȖ%��}�ٴ�Kı/����2kZ���W.h�r%�bX�g�w6������5Q,K�������bX�'���ٴ�Kı=�{�iȖ�/B�>O�ݰ>l6QQ�gy���D�,K���bX�'���ͧ"X�Y.Dȟ~���ӑ,K���w��r%�bX����{�:5�fkZ��m9ı,O3߻�ND�,K���6��bX�'���ݧ"X��z��P �R��?�*�L�z��&(����s����OW�z�z}�}��5�Зeͧ"X�%��{�ND�,K���"����O"X�%�����iȖ%�by����r%�bX����32[.��z/]Sm�K��FU��1ٵ�����\M0���ؤ�lB�F�)��y��Kı<�_v�9ı,O��xm9ı,O3߻��Y�L�bX����6��bX�'����C2kR�e֌�˭]�"X�%����NC�O�2�j%��w��m9ı,O����6��bX�'���ݧ" �L�bw���j��j�fkFӑ,K��>���r%�bX�����Kı<�_v�9ı,N����r%�bX���i�Xz�3��]�OW�zwIz0�"�����r%�bX�����ND�,K���6��bX�'������z�z�����j�����,K���}۴�Kİ�'���@?����i�Kı>���ͧ"X�%��~�fӑ,KΞI'�w^�,������E5�Bb�8�[p m�mz�k�k%anE��+����t	�����pR�:(��� �`��]�Mӷ��e�YM]��P+i�uR�W]���P�mږ(1�u	km�6�Y[��a	��bו�몮j��M�i�n3q)��B�V��\Z\��E�e����e��%р��]�F�[j�J.�3��˧�ݗ�qkK�G�:��S�s�l��\�n���&K�X�
�6�	\��PD�.u�����j���Зd��Mla����O�>ޅ�^������ND�,K����ӑ,K��o�iȖ%�by���r%�bX��t�̽��34K�6��bX�'���ͧ!�*���b���� �j%������ND�,K�����r%�bX�����r%�bX�}��UM��aq��нн>~����r%�bX�{��v��c���?}��6��bX�%����ӑ,K�~���ϕD
m��:z�н��$X�Y$bAr'�o��ӑ,K���p�r%�bX��~�bX�'}�}�ND�,K߻�9ɭK)�Z3S.�v��bX�'}��6��bX���~��m<�bX�'﻿�iȖ%�by���r%�bX�{��d���rL����go:I�^��s��3�IM
�*6f�fMJKM��$$ �Y`��>'��I]I�le�g�?/B�/B%����ӑ,K��~��"X�%����a���șı?~��ND��z���-��a�4�(er�t�zX�%����ͧ!_�"+��>D6�'"X�f��m9ı,O{�xm9ı,K�w[NDS��B�1'N��סz��`�֫A�-�"X�%��}�ٴ�Kı;߻�iȖ%�b_=���r%�bX�����z�н��>[���Ჺ�볼�Ȗ%�ʐ?����'����M�"X�%�~���m9ı,N���m9ı,O3߻�ND�,K�O�ٗ�#�Y&f�sFӑ,Kľ{�u��Kı;߷ٴ�Kı<�~�m9ı,N����r%�bX��wy��K�/�5[vڒ�t��2�ݡڰ����,�R��[kun5�S�﷭�IoI����0�SR�e�k[O"X�%���w�m9ı,O3߻�ND�,K���6��bX�%�߻��"X�%��I����f�ն\˙���Kı<Ͼ�m9ı,N����r%�bX�Ͼ�bX�'{��6���B ��L���Ͽf�u�ғ3j�Ξ�B�"X��w��"X�%�|���iȖ4^HOY�T�m��ѭ�y��.�Nl)X���_=�CЪj��82C�B�!Ǉ=&��||5��k	\0i�{_���HR�X��@�U�XD�Ri����j�؏���6,�BtH"2�P�)�(iKXMh��[dM5�⑨�.����&�xy5���LL<��M^U�|�����S�8w6�ӬŇ7�4!#�V���&"�a�H�"RR|�'4��6��C�,��$'�ǁP��e&#$!v�ir��KF�L�̄`؄����WJ�
�#�+�)�� ��'P�@6�hA��(��	���Z�T����)��%��|�&ӑ,K��>����Kı<���|J��h�˲�:z�н������Kı;߷ٴ�Kı<Ͼ�m9ı_�$�D����6��gB�/O�~Z},��)�������D�,N���m9ı,?�c�w��i�Kı?~��ND�,K����ӑ,K��!���&~��r�sY$�fp��,�,�%o.�u۩����hKf"]�gM�h]�=j��2�]?/B�/B������ND�,K���6��bX�%�ﻭ���"dK�����6��b[н��0O�+��
�:z��ı;߻�i���,K߻�[ND�,K�����r%�bX�g~�m9ı,K�>;f^莍a��\Ѵ�Kı/���m9ı,N���m9��"�L��~���r%�bX��{�_�N2q���̭w�%9H�)̹�kiȖ%�bw�o�iȖ%�by�����Kı;߻�iȖ%���0^;U_U���5���ki�нн?~�y(o�6)��|��%�bX�g~�m9ı,� ����O"X�%�{�kiȖ%�bw�o�iȖ%�by�Ӽ�ɚ�m��5ۢ��B�l�b�ht��%�;�mrYf[�\Li�fV��͙���н,K���6��bX�%�߻��"X�%����ͧ"X�%��w��ӑ,B�/O��~n>%Lmtler�:z��ı/���m9 ?A	"dK�����r%�bX����ͧ"X�%����ND�,K��K��\�Yn��]k[ND�,K��}�ND�,K���ݧ"X��ș�����Kı/��[ND�,K���f[�MkR�Zh��M�"X�~P ��Q?����iȖ%�b~���Kı/}���r%�bX�����r%�bX��m��|��]TTSΞ�B�/B����xm9ı,?�X���[O"X�%���w�m9ı,N���v��bX�&Ӂ9,��0��߳��y�$��p��Wv���Tu[��^���Q
U�$B۔S]��`m�m�6� -�Ŗ-ELmf�ш���s��,�k)��:U5x���6��6�V�ڔ��4��c9�ea�ۢ��7���]FRjjC�X���q�lh��#fJ�a�@eεæ���nͲ�V;[��z��z�5�:Z�M��_T͔��Т,2߲~��>�$��C���*�iN�Z��c�A�`G<��A��b͇M6E�mƚ�a�'^����L��M�K�6�D�,K�w���r%�bX�����r%�bX��_v�?�	�L��'wo~T����N2q�a����4�E��kZ�ӑ,K��~�fӐ�r&D�?}���ND�,K�����Kı/}���r*ؖ%��{)�L�˙t[e̹��ND�,K���ݧ"X�%����ND�,K�߻��"X�%����ͧ"X�%��~;��+JK�`��Ξ�B�/B�����S��Kı/}���r%�bX�����r%�`'�$2'���iȖ%�b{�M�j�\�SP�k5�iȖ%�b^��u��Kı;߷ٴ�Kı;���r%�bX�����K����=��Zas.�,Te���4R��Х��]L7B�jP��P�m��b ,مڤ���fk[ND�,K��}�ND�,K���ݧ"X�%�����REc}���%����[ND�,�^�����u��B1˼���/B���u�nӐ��+�$H�'�O�;���&�o��"X�%�}���r%�bX�����r%�bX����O�(�r�<���/B�/O���6��bX�%�w[ND��)?�� ��j'�~�ͧ"X�%���~��ND�,K�O�ٗ�#�XfjK�6��bX�%��w[ND�,K���ͧ"X�%����nӑ,K���w�Ξ�B�/B����>_N����ֶ��bX�'�߻�ND�,K�H)�IO�����{ı,O����6��bX�%��w[ND�,K���-=MlHѳB�`b�2���65���Q4`�ғ1��T+aCD��%#-��a�ə��r%�bX�{���9ı,O����r%�bX��~�l?��L�bX��߿fӑ,K�����93ZԲ�sP�[sWiȖ%�b}���Ӑ�P?�	���bw?�fӑ,K�����ٴ�Kı>�]��r%�bX�~��n>%LhF�Y�OW�z�z~�~�m9ı,O���m9����ҕ�-����X[F��@�M������Ț��Z���Kı;����Kı<�����f�.j��k6��bX)�E�Dȝ����ӑ,K������9ı,O����r%�bX��~�m9ı���_{εZ6�o�=^��^�'�뽻ND�,K���6��bX�'�߻�ND�,K��}�ND�,B�������أnNu�\?�1<��x�\\��1�c,3
�W9�6�f�4���.����N�t�,��Ie��=[��Q�1q��>�bX�'����6��bX�'�߻�ND�,K��}�ND�,K�u�ݳ��^��^���{�
�,c�ͻ3�9ı,Os�w6��bX�'���6��bX�'�뽻ND�,K���6��� �b�"X�{�~�N���	\�Ξ�B�/B�����6��bX�'�뽻ND�,K���6��bX�'��ݻND�,Kϻ)�,�̺-�������K��  dN��߮ӑ,K���߸m9ı,O{��v��bX]�'��c�4M)���I���L6H�tK,P�)�	G ��!����W >~P6h�]��L��d�'}���x�tLH楹���Kı>�{ͧ"X�%���#`�����<�bX�'~���Kı>�]��r%�c�߿�ώ�6�4�L刨Z^g���B�k%s��.�4[�!cۅ�q�3WZ�ӑ,K�����iȖ%�b}��iȖ%�b}�۰�U�DȖ%��߿siȖ%�b{�����3���K��k5v��bX�'���6���DV$D �\��,N��߮ӑ,K���߹��Kı=���r$�$Oz}d�&d�.Ys4��H&\n�&@�+��eBK�&Bq�����ӑ,K�����6��bX�%��o���Zmq�Ξ�B�/����Uȝ����ND�,K�����Kı>�wٴ�Kı>�]��z�н��Os�Qe�tٴϝ=D�,K���ݧ"X�%��~�fӑ,K���w�iȖ%�b}߻ͧ"X�%�SBEq�X%��H�Ha BHd��HKxЅDB
&z�f� -��׭�d�nu�NR#����b��ܶ[�6�r�M�o�� �mj�Jl�;Gm؅��Թ�&�)�-����T55��[6!��$�q�:K��5i�N���eٖ�v�4���v��s݋�h݉tYl\�1q�3\�5�xe�1�Л..������%�l�i5�5;�2ܥDc��+3	��Y����Ro4��o6	����T��iu��\�8ܠ�5�rm ^rĚ!l�3�q�>H$dPi���!��kT�E՗Z��}ı,O����6��bX�'�뽻ND�,K���ND�,K���ݧ"X�%��ݗd�d�e�-����M�"X�%����nӑ,K���w�ӑ,K�����iȖ%�b�r��_�^P�d�.�N�ߦGɈ��R���r%�bX����6��bX�'��ݻND��(D��duQ?~���r%�bX������Kı<��7L�۩�
jj�m9ĳ������Kı;���6��bX�'�뽻ND�,K���OW�z�z~{��z������bX�'��}�ND�,K�# ��~���i�Kı;���m9ı,O{��v��bX�%��%�ce�9�L��m���F%�2͔a�vX��]F\a�.!�ciCv�V�D�[�OW�ı>�]��r%�bX�w���r%�bX��_v�?��DȖ%����龞�B�/B�=���؟j5��W6��bX�'���6��1�X'��!�<W��=FX�R��%���w��r%�bX����M�"X�#���u�ᗡ�@��O�>�r^e
Tᙩ.h�r%�bX�~�]�"X�%��~�fӑ, C"dN��߮ӑ,K�����m9ı,O{�w�C.Y�R�V]kWiȖ%���0����~��m9ı,O�����r%�bX�����Kı=���r%�bX����,�̺%�������Kı>�]��r%�bX�����Kı=���r%�bX�����rt/B�/O���m�k�C�E�벶B���V-%�h�-b�gMuu��� ` ��e[�C'�=^��^���翞��r%�bX��_v�9ı,N���l?�W�� �5ı?w_��l�z�z���K�6��B6i\���Kı=���r%�bX�����r%�bX�{���9ı,N����r'�S"X������3���KsT�f�ӑ,K�����6��bX�'�뽻ND���C����h��T�+B�r� p
2l7�Rkn��Κ�AMݘ 6���=A�cO�r'�}��"X�%�����m9ı,K��}�oY5�Ku���֦ӑ,K��;��ӑ,K��~��"X�%��}�siȖ%�bw�o�iȖ%�b_zI�e;5u5.a�j�f�iȖ%�bw�w�ӑ,K��?�	����f�ؖ%�b~���r%�bX�g{��r%�gB���'O�~O��m���V� �eI{v�,����4�s����Y�p�m��f�5�-�1��hѢ��.h�yı,N�{�6��bX�'{��6��bX�'���6��bX�'{�xm9ı,O~�*� ��t�z�z�Ϟ��|���A�DȖ'�����r%�bX��w��"X�%��}�siȟ�����"��j%����vI�O�ˢ[)����ND�,K����ͧ"X�%����ͧ"X�%��}�siȖ%�bw�o�iȖ%�b}��ݽ֥��kZ�ɫ.k6��bX�'{��6��bX�'���ͧ"X�%����ͧ"X���:��x��M�?���L��߳iȖ%�bw��n����˅5&�56��bX�'���ͧ"X�%��{���6�D�,K����m9ı,O���6��bX�'���d�[�`Mn���]�e�bR��e$�nb��"D�j�U�յ�k����2d�󧨖%�b}߷ٴ�Kı<�����Kı>����r%�bX�g�w6��н���_{εZ
kL�Ξ�X�%��w�ͧ"��\��,N���M�"X�%���fӑ,K���ҙ~8��N2{��Be�x�3�5�ͧ"X�%��~�fӑ,K��>����K�"w�w�m9ı,Os��ٴ�Kı/��~;���4R�%֦ӑ,K?�@���fӑ,K������r%�bX�g{��r%�bX�w��m9ı,O~�<�ٌU 0A˼���/B�/O>�fӑ,K��;��ӑ,K���o�iȖ%�b}�}��r%�bX�>MC�~_@۠�z<շ�G*�+�8CY�R�y�{4q߮m�xIO5CZ5���1$!$LON�i�o�8��#B$ ��Bf���@#���8ksD�
2�Ö0dF"�8ʺ|ʦw
2M]|���xC@l�򸛤���Bo��403���v����R���L<�M��!<Xl�}�a��ተ8'}I5hW��d����S��' Kk�/w^���� ���� f
�6���:=� Ѱ����^����` [v��h   @ l �     �   � ��m�� pm�@8 ���!  � �����I{-n�&5�ՍY3J��M�2l:ǆ(iev��Nl�eSVΉl��#�����m���6i�).���Ap�l��9m#h�8	 ��    �   �����     � -��          p      N$[n���4� ��үku�۔ơ5�"/k�]�X볊iP"e�*���[�� AUrR�U%�\a�T�ڀ��)I��6[���6P��X�cҍF�:m�j�  H H[E�Nm� R���"�,��Sv���fQٓ2l[Z3h�u]r]31�Mئ�YB,N1,J���Kr�M�G7�s�,\��	nڰ��u�-����e������$�Y���5�h�,�#4�f����&��ecI�rDB`e���6H��6�:R�ܓ:�h�n��.&M�����1�I�H/R.\-�鶵�vچ�a�q f��	����K�F15�p�Q�Yj�j8��[�r�T�m�J�A6)Pfk'Q*,�˛ӣ�t��N��{m{H�.�&�����a��\��1���:Xh)�%U�R
�R�Ɛf�6����U�le�m��fd1�Y�f5�*���"b�\,Xԧjj�"�@�5�m6;U�jj�]�H�k�C���G[t�M��E.��ۑX��E0ִ����/!I���.î��ک���C7e��WQ��IF/L�[	���	5:[��ָ� ���A��0�`6�ӰA��x��&-�F���D]ڴ����c[�m��"���tٲ�Y�s:E���;�q͵786)h�dH84��S0�a3�Lҗe�LhXL��Qm���k�k �efiU�Z��E3v���0�3z��r[�tpD��D7A�6
TC�8!��?)�<@���B��CXz
�'��|=&}��n�v��6���ڢ�����KM.YfJ��(��a�v��eQEcl�U� lݮ��!��6�"�m0SQWEuea.�c���:] @�٬�!������Թ%�6��5C\�(��\�P�Lкl[��t���J�����`�L�l0�m�ҥ�D�t�M��Lm�FpѮ�ً�.�t�q���P�nu�*��M�=�:O��I��ڄ��M|�k�m�	p��̫eM�3i��l������<�R�v)(]F[�]��l�\�����bX�'�߻�ND�,K���ͧ"X�%��}�s`��șı;���6��bX�'{��V�m��Jgy���^��^��{���r%�bX�g�w6��bX�'��}�ND�,K��{�ND���,k7�-S�H6�L����|r��G)	��fӑ,K���o�iȖ"�Dr&D�?~��ND�,K����iȖ0��������.B�L��t�z,K���ͧ"X�%��w�ͧ"X�%��~�fӑ,K��>����K:�z���`�֫AMi�����T�,O3��m9ı,O���6��bX�'�k�ݧ"X�%��~�fӑ,�^����O�~�-�m��á1��@WX�^�%�c��*�r���j[-ڤ%��6Ά]� ��byj�6������^��^�?w�ӑ,K���}۴�Kı=����"�șı=�߿fӑ,Kz����'��V.̢�:z�Љb}����rl8HՊ�֌hR({	��QC� ���<��K5��6��bX�'s�~ͧ"X�%����fӐFı,O~����@`���OW�z�z~~����r%�bX�g{��r%�bX�{��6��bX�'�k�ݧ"X�%��{.�2��ˢJS&�Z6��bX�'���6��bX�'���ͧ"X�%�����iȖ%��dO~���"X�%�>{���5��[�;Ξ�B�/B'���ͧ"X�%���}�v�D�,K߻��ӑ,K��;��ӑ,�^������奷;mlm�D\ a���&�u=%�f-�$�U%4-{�y��e��5nfJd��33SiȖ%�b}����r%�bX�{�xm9ı,O3��m9ı,O=��6��bX�'�����S5�fL�ɬ��r%�bX�{�xm9,K��;��ӑ,K��߻�iȖ%�b}����r'�S"X���݃�Z�&���OW�z�z~�~�"X�%��w�ӑ,}p?%R� �V�KT�)�"n'w���ND�,K�{��ӑ,Kľ����_�RQ����н���Mz~����"X�%��뿮ӑ,K��߻�iȖ%��  IQ>����m9:�z������G<�WfS3Ξ�X�%�����iȖ%�by����Kı<�����Kı<����rt/B�/O��߾��pkg�ʰ�����\Z�̩��BkL\��ybm)X��kun5�P[�$�*��S�O�нн?}��ʙ~ϟwb���t��a��ݍ�3�
P4�R��L�J�>[�����$w6x�7^�Xw6����1e3RM�!Pi8���K1�=�W).���������DT��m��)Cn���2s^���iP�3"��$ə�3�C���o���rO���~����f����`}�۫�+����?��l�`}�5X�A�H�i� ��"Tid�4�Zܗm���CM�M�qKa��JiCi�л`xA)6��`|�5�w&�u�y$!7��Ԩ5�:9ȗN�f�������@{�T���1 |a��(�"���B��3�5Xw6���h�~ފ�g�������䉷)4)"�>�mՁ���`}ܚXs��ܛ�`g�*�h<ڔ
�29*���-�{�r�� >�ʭ�0ѐ,!	�cq���|f�"�������@�M�X�)2X���_[o�V.�bAʪ�P��m2�z��oF�Wi3���a,أ���<3If�e.�6�WͶm� [@&uc6��r��1��
6b�İm�2:�2�A�f�	��泴��k#��<�YA�K�\��okcGF�k3ie9fƮ�]�ʚ�*m�Kuu��[[6�&�w�H��H�"��8�6�3���m0$�V�\L�f��Cc1t̵*�j��5Q�4�sW�I;���~N��C_^�-� -[����ٰ�XZ\�5G#6�ͤ��q6���Ye��O������]3�n9�6�X��O��}�Z���9h%�u6�L�.��h����@{�T���-���+�Č�������t���8��J���x�y��&�Flo=��@j5���$�Si8��y���㖀}�Z�E� �C˺˘n�]ʙ�w�z��Ǡ<�7�^fd˷�y����l�>ך��sQ�T�
�P�c��M�uX�-��0F��-5c��t��A�CMc4&1��9Ȣ"�8���Vٻl�>ך���V��6(�h�6�<8�2��̨*��켛&�L��i8>!�*H4�h�8L�4 P �8�P�a�<<-����F�`T=S�g�Ͻ��o�x���^e��2�D�:���y@��!@_F���^=fN��|��}a`ohj��A$�q�FԖ�}�Z�9hG =1�@zK"�� �R�N+:�U��_�U\��������3�5X�[bi�+vX�
����U�4)E����.ڔ-s�0,��� 6����;9<������Lr��K@>�- zY3.����T�7��^j�7�uXך���
乙�Q���u�L�w�3.��dw=E��(ju�0��2@[El�`@�#c �Պ@�_5�;�ɹ'��~��t��s���8�=�W*���+���@zc���d��|�ܼ��ݸ���'���>��Ǡ;ɐ� L�fM}[�������@y�����G孉6hQ̻\�V��in���F
�]3L[,X�fx��"mF[�]�ZBl:��w�|���U��y�ܮW9�n����P�R��D�q�FԊ�޽�W��發�L��5Q��y�ޠ�?\Y _؈�%H6���ӊ����V�m�����`o^�;��Z�u�����h�@���1;$�ڕ���O�4��O(��)�]�+ ����_�R	H��n���1;$��r��������~�6��XE���m��2�$��J��b+��R]���a{i�]6�Z�J�$*[���?����@F��9��["�r(���Ru��?ʪ���D���oE�d�@_׏S*!2D��L$���Ͱ�>[����,��Vf���&ԠT�n@�?>^E�d�@_�x��&B��t,�C�K��&�s��G`ovh�}�Z7 =q�@�}��KYY�fH�Y�l	���R�-�Y'ے��I��דW�3vA
@��Ȫ��ͮ�nͶ h5+�v��u��L1�e�N�n��.�D�k	eUtd-�M)u(�m-�dqW�����aܖV��R�[{j4���m����*k�jfZ�c-lMd��K�!�N��7���n]���ؖޝ/#�đ��v�0+K$�"�Cf��Z�g~I'+��;j]��*S8X
����4�Z�b#5��1�h1��h`��;jvG[�o�~���h�@���1:l��I]A���U�73l/���W)��w������qx��ɒN���û�
A):M��:�|���,��s6��;�,kXʉ�$Bq��N�Ǡ2�((9y��
.wz(ƞ��(�"��85!`}�5X� @zۘ��6	r�u�3.�7+CA�(ە�[���������A�Nn���%ms�5JE$Q	�$���+s6����1:lx�����,��ڒ�.f�&䜾��o��"D��(IHő��Č	����_��d���y�~��~ݞ(��
�$��b!:}�%�"&%�����9�@F�[swQl�b�0m���6i`nf�P=�E��BaGg~���~xw�#�����,������w��=��,�f���^�#���UQ�A]�j�Pt�b2�Ɔq�D�&�u�k�Ȅ�� 	�JT��S���Ż�`ow`��n @%X�,�i[y��q�b�ϲp��Bf�}��z������UT�i�פQ�DJ�87�(�7b�˼����i$$��̐»F%OC���FzS���&x�|z�=tp8|I$IS�	�P�8s��$�=�_�����>>|�R>�E�Jr�$q}JE`<-!@0�0a!'�#H�)Xp�i���%
���}��a���!!]y(�6�@�H�����Ag�j���ۅ4z��;`4���G����6��6B$d4���
 :H|��=�@�	�����8s��*m>~�}���Զi�pl�l�g8��t�`j!�p�-�8x񙏬(ec�E�lk*x��	��8��{��㨺"�ӣ<�����m��8E8"�@pE�)�<�
�"x��!���"b�6�4���W����ƒG��� �)>8�T"">�x�T=U�@>9�ֹ���K;���(H�r���#�2�((�w�@~̜(9�30��Qs����ߒ��BmJI��噮��6[s��������U��̡�`��Qp����\�ЋoMy[�lv�V�Gi�L��������u˽�������n @zۘ��K5V�q�)�&��噮��������z��/w��ϲp�>�w��yw�faY����@�<���@z�5�ڵ���IH$�I��f��d�@~{�����C&K��{�������_�eD�RNK{�D����?g��'���@{��m�5�j�	�UmU����!V�&���33,�,�-V�g��3�O���"8Vyc��R~ �� #q �sP�� �˺�I�w�@L��b�˼��d����M2��=���Ƞ>�w���6���r�}��������fk�73l,��-�&�s���X�N�Ƞ2�((9��a	�g7�����������lp�>ך�� 󘀝6���i2���<"m�Zf�����
�r�d�aP1�m�T�^����u��14
L��m]���m)�y���[�(j̛nVa�v�cG���mv���m�/�� �2Y�����[rY`Mk3�R��P�9azÃ.],�Gc[4������ș%q53Ŧ�ZV �TT�k�v��h�(�
2��ہf,v�k�2��k�1��-Sk�"�i�I�8�9$vl�u�-ۥ�Ϊ�-LT�[�e�f�6���~�(�������3XZd&R]]I��e�Jܬ6RBT��R��R:���[�l����R�Ce1Ȱ�m�����������^j��kImB��I�N�p��@N��9h�@��_j�
�ESa��^i� ��$�?o����n @;�1 �u7n9ȉQG�,��s6�����`ovi`osR��	NPRR+.��d�y/&d�����������W�Լ�iP�n��'țm"˅��e[*lI����]L	[�&�v�mt�0G��6��Ԓ3�5f��ݚXk�^���|�������JT��nG9$��>��}7
�J)��"�:a�@��T&���v�I�;��ܓ�w�Z�o37�HBd	3L��r]G���("^ ""J=����I���>���`fbQS��BRhl�9�L�����1�6(�'
>�Ǡ�kIV�))�J�#,Y��ꤼ��0&���|dw=y�RP�/n�m�0.v�QX�
�D�]	vX�5 �]�pZ��4͇$ژΆ���R��[Vݛ�	�`���Z7~����� 5V�H�� �q��z�U��T��͠�5�6(�'
ԓ/%�L�Oo��E��Br������������ř�sJM�)*�%Z�PS�Ns��j���r���4�;�uX�JP=i&�
T�n@����qk��=��,��UW�}�X��)R�$I��.�m:ld����2K@|���=��|��q���!p�����&�u���3]���Еꮣ��Yq?��t�Ζ���j��8�q6�`����73l,Y����U|������Ԣ���BR!D2�]�jfd�k��P{:P�uXڵ���IH$�	�V�f=�d�G���&��@owE+ 锱�j 8�"R+{�K�3��̊T��t2I:�:fN��*�+�<�v*��r��85 ��$�9-R[��� 9w���,*f�n�RYWZK��֚��	���-�Y�F;rJkun5�&�:}�[�z�%�$���o�~WV��U��٥��y���jR��I6�R�ܑJ�>��M��9hrZ������H�r9��XݚXך��꺰>ך�����!��mA�m���� ���z7��P�/��̟/kJ=�EO�҄�:l�r+�����9h�`�}�Z}��U�R̽6��՜��ۀ�l�������p�X��,�X����JD��EV�:ޫh 6��K��7�fE�镣�fƺ��GU)kփ0,vR��CK�F�khJ U��j�l��]�-yF���R7��Q����kCv8٠�j�E.��!�3�ZQ�����U���a[�!km��ј�qR͒�f�f�6�g.�2Ո�5t�6N�d�:շ ZSΖ�X�
�[�p9�f��6k�æ�f֖�Y����i���6��0g�]�Ҡ/�(�/̒�>���zT��y�~D�"NJ�3�4�3��9�j��*@K��v�6�C77t����@s�� =T�}6njJ���I� �b�X��u`~��T�����7+y��w���6� M���ͺ�?ʮnz�|��+������� q����T��Z٥� V��;j���Ŵ�2gm4l��a(K��)�m�9nwf�c�Vsu]{���wޞ,�j"��lmC2L��ܓ�s߮�"�M��EX��Q� 
���5?o���`{OŁ�٥���QS��BR6q���ݶXn�,��W���`n���I,�))�T�N2��vi`_�8Pqx��̈���
 �w}�s� 8��wf�c�Vsv�`}�4�>[���
��AR����i���9��F܍ ��͇M6J��k�1��y$QʐrA�1���l�>ݚeWXg����IU��I9QRM��hol�z��x��}�\�y��M�;��DH8<D��{�‿�p�W���@�L�&$Q�W�➈�9w���I�}���f��-�6㜍�;�K1��̨(<�3?ٵ���r]F�& �y""$�>��z̗�c7��>��������7���M: ܔܠT�A5�)Vh�kC5��9��\�Fi��q�t�*B����n�,�f�wf�q� �V���))�T�Op@y͂���U��� ����+L��#Q q�H�p�;ݚX��z52d��̘Jgw�NPޟ:��r��jB��<�`w����sߵ�ܞ5a�8�)	S0hY�)1
�"}�-��z��[�ē�RM�E`w����� ;����WI�j�)#]�s.�!�����4b��[���J���5�$^�2*��4��$ۃL#��>͘P}������y2�r��r�����J��!N9��p�;ݚXǚ��+s`��f�J���3/L�����@w8�@y͂���o�~�&��t*�!W7�������+
s�z����@~��Td�3�ei@���B�r�qSMӕ`}�4�>n*@s{����UW_W�}E^������O����7�J5 B!$f@c�B���k���4BBD�ɣL�͘I�8��o@������B�%jk���Xxi���F2CMʭ�$d�L�H9�)@k�*��C �bMV�Q��	�p:L#3F`�k�S5�LMb�p�*�a��`�vUպ�Đ�F'��h���da6���8Pexp�*>a���oFW� ���"B)�*ECjj�z^���zw����0�n�Tr��ܛQ=�q�٪���u���]�L/2� ��    H m�      �   h H�����	 ��h-�  �` l:X�[�[�[l���El4uFa�*�&�1�6γKGm�4�;�7TDv 2���vۙ�=SC2�p��ά7�m�;��angEۖY��� 8h     �`  p?O��I�[B@     hH �J $         �      �l�hp��@��Y0�KdF̩����i1��^�j�o,u�m�[�;E-U��KCZ�W0aGv-r[�ͱf�)K���e٤z�.�I6�6mڮ�gm�k�   [D�pl6�+T�[��h�l�&��(�;]6ٶkX�3��0��5�������n��VU��I��W��%�d�)v��M6�FX˥�����B�,pbY����3�(�_&��3bu��[�P.�4�vIe�U.�%J^�m��y||��:�0CJZ�3
��ڨ���J�%������HW�M����6t�N�GIɯ[�@�!z�������3���ɛ�[fۤV�j^��5��X�P�4��-�%F���^lV��R�GBՀ����`��t-u���tt�l֍�4���\�6�Fa���g�E�6�hֱ̤�bR�!�E)h��idԢ�Kn�fR�f֬ѭu������0��cH�j��IN+ZWD�kX.t��kf��`�0�Hb�[� r�+t*]kJ�$�SK�[%��p�YjEv�s��\��Hr��\'&�*Љ��u��ZŸ�m2���fip�.��A%s���:�i6�rI���Ki.XcT�l,4�ڵ���Kkv.x�c+ZvRX�ԋ��N])eu�����ڮ�v���Vi[;M���'X��\Fe�M
�Mu��f�&ذI�+�䛍f���4b���Q6'��UP6 uM�q���uW��D}@�#C��\S�4D~@�| �>�������t�-�� �	�nU�ij���5��t��j���[$Š�l�u\6ٶ�m ��0k'5�f��ͦfͣ�n�[	�it��ס�I�_��t,/��F�;�-���Y��][�̤�A����Bmn���Lf�@��M�0Ò���mZ�l0��GV�Fm�ɮh�i]�,˷l�%@".�ԫ���U�3�
0�nt�U��Y��;��$�?:N�:o?=~Ers�"���m��x[v.b��aʔJ�V���b�L���$�ݡ��pT���"E��{�Vs&�ٛh�>͚X���dQʐrA7*��d����(��z��/zx�>��Tس�=Aē�RM����3mٳK��u`w2i`}�J5�1�6���,ד���R�>��(9���{�(�D�O�$�<LKL<D��yJ��fd�9��t���9�@�s0���ƕ)�,C��:ʴt�k�k6&1b�6jB�.#���v�Vym���}� �w����p��%���6������S�Hp��H�`gsm�\�H�6i@}����/��%�7���ߔ�f�qSm�U���?w6���<�`gsK� 锱�j 8�n�?f�y��^S��3��ZP��^�G9 8�r;��K;�h�>͚X[��X�Ԓ�D�(�uj�@�ݺk���m��#R�D�Jsvu��\��}���u���I9$�:�߭�6�� 9���.�2^a�fٙfV�n9�@;�b�� �2����#}�JT��Dӎr4�,^���{�8�����0怉��ж�`G�	M��W4�X�a��ӎ���b����X�JE ⏢r�U��*�G�m�w&��Z��#��̼�3�(���P����i`b��`}���9N�!�B�#�w�PPd��ͭ?���@}w8P[�߲���w���]�j�!��L�Z��!���"k� 0ݖ�qeթ �8l�f3J�I�Xf�,��Vs&���W��u����e�i�^i� ��H�p@>�-��8�@y͂�q��(�$�rE`w2i`f��,�f����Xjpq$�T�bݴ�-s`���Z��U>�UP2`V��q�i�WH�q���)P�A$����> uC�����O���L�Wׯ@n뼄y��%��"SrٳK��7��3^�Xnk�[����6چ��M�\.�+x��:�"�\E(쵂�,��ͫ#�s���5"R52q�F���{�Xǚ�75��٥��kT�Dq��R))��y��3s\�>͚Xך��UU$w�P^NS�Hp��E"�����٥����������i%��IM�J�W��������@I��:e-���(��H�p�7�uXǘ�y�@~��(�$�	��[ҝ!�K����.�K�&��r�f� -��׭�d�n\����<D�i��r�,��r�mpz�� -��%�&햑9ykq
.�*�!���hҚ�ܘ�V��И���f�,��gC4����m%8�$6A���f��[f�Y�CY��`�lغ-��ttĺ��kuy�WY��f�v�α�� �X�f�o�3�㉯SO)�F�V�3�.-���&D��]�j㻺G]*�Lk�.��6ʨ
��Kx�4x�ff*�r^ł�?�-�%�V�����%����}OJ9�nr��=�~�o�����`}�4�Nr�_ �?yX����ē�RM�E`��_���T����`{����VsR��lLq4���sP�`���Z�r�n�Z�>4���1-/P{ɘ�򻞀���|�$�>�֔�Ǒjv�ґH8�ǚ�s�[��>������uXw*h $t�2����U��Y�7*g2��� �*Gb�-�{ZV�Rk�(��Q�HS"�Xf-��f��{���y���^���P䦜�N\�ַ$�ϵ���1'`@`'�T�%�&f^�L�ٽy��{��.��l�Rݍ�D���{��ˋǣ��$�fc��{:P��Y2��H9"NH�ǚ�3�{�Kܪ��OyX�i�
��Iȩ&�%���&���okO�}q��\^=��Z�bT:�]'țmR�Ԃ�̫b$�I�3]���-�y4�6�M�Ґ�ہ��&037r�P����-9h�{,ܨ�Ky�q�Dۅ��^�2�����&�ϲp�I���IL�˞J��ԡ�R)'�����V��e��HH�I$@H�H1p6;>�+�_u�����}w����uN�����31l�7�K@{��9hL�ww4�wk3%*q8��7�uXܮWs���=�|�3��U\��h�M)n��Tu����\���R�s���jKm�F��֘Ά>���9J�K�CD	D�R,}�?�./�.��|�~pۍנ5��e�%IC�H�r��V��e��{����4�7k@��r*I�H���	�%�=�`����]��[�C�#��D�<��ɼɼ�
}���3}>(��(��3�C�����L�B$$��(|"�����9ʟ-��|�H{�3�Ld����� ��@N�-�ﾪ�>Z[�mln*s���	mh]n�p��$5��z9VQl��,���ka�h(���x�o� 6�jvIht� >�PZ��Q�ȩ�8Xf-����^H�;#��Ξ(��(���%Jm�T�qI`o^�>��,̚X�� 锷cCD	D�R+�6�� ����Z]2V��i�QD���72i`}��vIhs� z�����^�yy������6��כ[U��[j��:�5���1�[�핚�M���Q�o�� � ����n����]�Sb �kX��7�%��V;)JP ۉm!k�Z[[l8B�]]�Av��Sc����6�іQ�CJLh�t�t����l�q03rś$�fƍ��1�`��y�-�!�դ`ں��e�4�1��iP�[�˙���u5��
�<�#�RwId��<��������LՎ�R[\�t�*h��Mc	���1�\Y�F;KX���Mfj��7���l��������V�ɥ���K�F�SK[L�PIv���*�I͞,n���k�UW+��T��Dӎr&�Vsg�7�@y㹈	�%�:S� ^mf:R)�p�����y�~v�������1Aju)�E:r.G!`}��bvIhs� #{�8��aiLatq6X�
�o4�s��;he�3�æ�u�-�����1b�eVm�M���.K��X�m�hݣ��fƆ�(�����KUG9ÔV@� *�$�!'� +Iګ��??���������w}�`}��W�����y�N���%����Ł�r��W8�w޺�;�<X�a�.$Ĝ��l������=h��*@{����(�me�̸�!	�Iz��R�97����|���`}܆�{��4�P���Q��V�, @Vk�������0�d�����e%
�D%9�q�('%Xw&�s&���j�>�۫�X�����)������礴����@}���:��"���$p�>�CU��}��ϸ���#��k��d��x�v0��RZOtFA�t��XB+�Z�z9�L�t�B!���hy��C�	�p���BT�$a㫐�4�63F��xrVх%#0$�1�u���l��B.z�I"M�"���J+*�����+3�?��К��SF�UOO���Mm8l2�ᥱ�X��끳T9�0Z'�z	��Mi�D�R���!��=7�!i��\d����M��8h���BA�+�Q�055���H�$Xp�4˷I�
n!���c�� �<صD8/�������>+�'�; � �'��v8�T@��U�A�^. �Ȧ�5�$&|��:P�<P�2��E/2��J�nXW9K��}Vsg���K��5Xr����"J(�rU��{7�@{���r*@s�0۩ĝ}����m��+��rNY�tʽ��	�*��bļi�f����jh]�-�>��(�\���̥��d���g�s��Ƙ��RI���5Xr*@{����(�me�̼+l�ʽ�m�"������zj�3r!-�$q������K���ɏAmI}䡯�2�JD)fE"<_T���|��w�rO=<�B�CN��A(�,�M,���P�7����Ԩ�\�@y���p|؈�i[�͘
������t����R�ap��-s
�R�6 � �M�Xe�U��9��@yȩ�{�UU�&���I/T"��r�6�"�>�۫�����d����W��s�H3h��CD�(�$Q�Vsg���K?s����}���~�u`b�6����#j97�@{���r*@{����j�LIȩ$ㅁ�r��v����4�32i`NW+�N���4��9R:��՜ź� i�b)�ţ��Į�K6+�ƀ�hK5�PUMvv�L���6� -��c-ڃm��0��+մ��)ܓ���|J0-%u�fsX�i����4��v�I/.ڗe��i�� v�+n�������)���n�bA�ݣ��.�lRg6�3)��v�ƴ�����IMV�Y,e�j�6tu+ ʦ�j�HǪ�
G$�+(�V�*�;�;Z3[5ݠ#.�!���Gk�V9�Ks4vriY���E��^��tp�S����0f�j~�>{������(��?����J�3zO=�t��愎9�rU��ri`fd����Vۻu�UČ�j����)�Q9(̝(�\��k$����Tד�����S��NGN(�`}܆��̥@~��
&�Q���/���ߔ˾�^���ff�h�*@{�� ܊�w!��Ż�"����R9�IQ[k]�-����)Ya�b$��R�]��35�����v�\�R4��J���f�Ձ�r��s����u`j�=^iF��)��kSrO}����R��1bPqG�|N��A&��N]���]XnmՁ�����r*I��T�1��2��2o�{�J���������䦖��R���������r*@y�%�$�e��M�������ݤ�9h�T���@wwn�������N�'���#��:ʴt�k�k6&1Z�s5� s���A&�Vf�Ձ�<�X�ۯ�]a�~����A~N�:���t�rU����6x��R��2�jD���M9 ���,��Vv��dIH2J�S�?G��Ձ�ɩX�F�hh�"���h��Z� =�h?�_U[��x�5V�4�bt��C�X��V��m��������E���a3�д`#�Uoi��b����Dv�X��2XD%�涤�Զ�&.R�g���˴I�@t�- ܊��?��Z�p�JS�$J��������#<��������&�~�W8��z!/rH�g�x�(��z/2��7�y�)����+����,��sj�CN��A&�H�T��{.�͂�N���/X%T�G�@�Z��ryX�-N�:���t�rU��ɷh����r*@����6���X��i	��lnh �D�&*Ss�W]c�p1A`�&6P����l��@G"���v�=(�rƉ)R6�`wj��W8��߿]X�O�Xǚ�U�kZQ�:JT�'{���R��v��Z�9���PbNEI6��s�so�X�|���v�R���U��Q����$P�TA3.���@y%�Id��|�u*���z�X�a�0�����޿��O��*F��8Ce� �T�Kf��M�cF�d��Ųr���Ӓ��An�)��6ݛl ��Y�-��sgnvݳ��CۮтkYD\VL6���ٸ�vآWfbio	P��hm�u�膰m%�,����M&	���6�b������\�&����5.\��*-��aR�λ;@����(.��������-�X�mJfݘ��mo�j5�*�����6چ�q�K��n6V�4Ky��_4u8��h\�R����))���53��PjE�<�~�`}��Vw&�`wj�>��ͫq:R)���f�Ձ�ɩXǚ���vw�R�DRr:q9*���Ԭ��V~�%���`w}������RR�
��J��UK����S�����w���y���s���ѻa EID����<�`}� <�˴���J2 ^^m���*�*YIo W`�{M32�H�Y����K��_֐��HU%F��_��]X7���{[s����e�������s����n�1@"�"ā X�"�≡�?��,͹‷��?}yJ�����	�#w4����3j��@s�-�qR�{��݈�8�s�E,?ʮ}Uo$��y?Z�$�@{���N��n!�JE �r;��`{�]��R�͞,��v�jh $m1���+6�nݽ:tB�������u�^mf�9NN�����?��O7���h��.�?-��7��h�@G�ZݒZ�����N%%)**J8+�ɥ���U��^�7h��F�i4FT�RQ��d�{�}w$���s�==b� P�B�*#-
*�eXUy� �#�!OU=TO�������3ri`j��Z�GI@��7���f=���}s����7�2J}߻�@o7�8�H�<L�w�y��3�Z��㖀�d��|��faw.�h_!���[.���ln��[I�6c��F6b�W�J�kcZJM.�h\ي��'���`���vIh	��ZG���N8��G{�K��)#���`m�-z�p�d���d�\��Q.C�)��,���V��j�;ܚXܚX��K]JT�I��ĤVܪ��M�+3g�{�KuTUN.s��B_�M������ј�I1SB�F`�+����8�Aj��UU_^>�>��6�ӉIJJ�����;ܚX�r��~>���`o^V�-���-���gK�V*��7[iWa�0jC.�ɷnR�MZJ�Zc:.ҫ��*RQ��`ori`}׺�����U�E�Xn�~,ʼ~��GI@��I�ј�䙝͸ů@]��@g�8V�&w3y�Ȧ+br$�R+�����6	�`��d������U���Ҳ�69QXz��U,Ϳ�g���a��Us��6��{b�B'nqH����\�@>��e伙f��>���?s�{7$�_�_��EEW��EEV�**��(��������آ���""����@�"�`*�,R���"���E�"�`��F"�", *(���AH",Q�"��",�"�`*X",�"�B�
�"��A�"�@�"�A�"�E��AA�"�(�",�"�B�`��(�",�"�(�`��@�"�� B�(�B�� �"�D 
��,@�F�F �@�"�@�"�@�"� �EF��H�� � �@���",D 
�T"�� �@H�, �@"��?�(����QQU��EEW����TUx
**��(���Ȣ���⊊��
**��(����EEW�EEW���e5�n� )O��!����}����'���:   �    )χ��  �CH���Elh$ 5)B�( 8x 	���(Q<��G���LhP�Z;Ra���pѯF�S���t(�,(P��w�� B��xz��^�}h�T����5�L �h�5Ѣ�]>��Ϯ}�2ɯO\ ��_iT���*��A&�٫uW}��]h���]u�]�{�]���=��9�ou�֡�}�>��trz������ ��5��M�}z�����-B�����h��w@�h�ـ ���s}x=q��4(p�+��:kC=w��� u����ӧF]��]:�tG)�t��]�a]:i�Zb�:t:>@    �!���J��  �`& EO��U�FM A�h  ت�=U&j h�  22   4�j��i)A�2 1 � 0��� � i�`��&�z&'�� �!*��      ؇����7���o
ٲ��QAh��C���PE�?�Q�`D�P[S��#���/�� ���p�_����N�����,����g�����������:��ѷzkݯi��i��X=�<�$G�N�PP]��i�"�4���MUAAx�@�Q�jp�fӮ�t�pa��l�&�0AP] Y�X���ߦ���٦>����ʨ(.���KM�����Y��Ѣi��]�æ��Ҫ���E>���4$�}�=l(6h�:�moR�b�I#L��u���ʾʝ�(�7�Gw7���7�HY���T�:�Β�EG[��HG���[�M�HH�	$^��A�	wʕ�M%T�K3P��|;�G���n�B񓐩EJ�vk�xo))��8��*F�!V³��%h���wmD��i"D�	$`@�J���X���|!�����˛���-�	g�%�5 �#M��@�62IT,�1	���m��ě��:|�4���&�F���-:��~Fy���4�JHB3�Xt �LNT
I�K��j��t�ht�1ၡ�����3d-�9ʪ&S7U�����٭��a�	�<2�I	�!@e:2�5�fP�������ƁE�rYpc�I�FH��Y��h�F��|��7��7�0�FbUU�[j4I!5�s�0��q�M�)�&,M�"xU��֤6cM$�Ta��/w^Ww��nL�^�A�_,�&���a
�
&��xM��F�Q)�^����E��!UC��	#D�Z��P�^W�d�l�::n+�m��M�ăE��3��Hj�TԄ����o�n����%�+.��D��a�B�E�2\-,r4\�q&�edz�;d
p#EƜ�:rlZ;P��=��<�OB6fJN�ɞ��w��fCP-!����n�^sv�!�g.W�3!P�e_Nj�B��,�1�fY���n��R@��"D��'>"k���H���D"� �	A/�j�wV$ j%�q�4&�Sn1�
	MْBNJ��O��#u�;\2<ʆ�U+e;�$��;����sZ�!�Q�[�4ũ0Ӫ��7�ȓ�z�o�K�.QX@�yƝɾ�b�W:dbԧ�$�w��D�҂�m�5 `J���a"�3���;	���J�C3d�$I��ԑ"���F�jT6��Ms�n9S��C�c�dnHF�Q�t�rq�vN�(d"B%����9�ߊy}5�Y����=*��+4H�lb�BHNh���HIJ�TY�G
�,���P��Het�8l�s4l�I$�p�J/Y'�Ӧ��]�*�0,m6M�v �nXw�8�����FJZ+KՃA��$kG�w��E�lz
)�k��R�\>BĪ��)X��$C��D��H\�A+$)��s����(�k���9�p�ܒM蹍|��޵�RꙪ�w��ݝ�����.��Uә�ƍo]8L��\kEx!��5	�W1���u�To:p&�A��	��cB��Ṗc(%H�,|�7���6p7t�ĕ$4m�Vg��rM����2��0��ץ�'�B=|U[#Z!4¥�mL���(�$�^�!7Ñ�(Ԋ��8�rh��n��(�6��5��e^CR�o	E��J
�h��gw$�n��h��zU�K�S���\JFvp�pγW�A���zw��_�	Hp�7�T�7n@��kr���v\�.�Y��U�d�q�DvcP!H�#I!tkN&�&�B6�D�6��dJ�M0(��a�C��qĜ�S����C�w�H:p��r�eC���些0�Rp��[��5�B�4LwY�I,����Fl7����i1�V�G�V���hQD��u�w�&�d��wxF��@���op��IUF��U�/�5�S�T8V�Jf�G:�|�����,���&'(���6��X@��5i`�j����8HR5p�*Y��G:�h���)�#��FB!�]��%VGD�Ԡ��Qn��c��$�9��vx�P���/5������05�Q���P�M����)��D��9����r�r�
5�P<d'8oY�g	f�'C)����#��0^�2G�#���;6�%I1a��F,<:�V��IZ�hL�ʜ+;ٜ��2����\w��eJ��\w���0+8�:y����ig)��·�:�P�K�	W��rl�(��I���m�B��$%I0��i˳��m5��nWt_��k5�4��3`@>8�.v����@�z�8N�����0���c�gͧ�z�S$�&\.������Ϧ�T�J��P�R�n��Rq%K墍�X&C�Z�	`�<��٠�*���{&y��ܺ�L2�&bm�j�Kx���ݰ�� �� q��l,�nP���	��f��m           ����      �                   �`          8 Ot<    �         �           p  � @     [@ [@ $    	m      �m�   -�   8                u�^�eTji�it*��:��)���K7K�$���s�~-UT�&�en�'b+T[��X�d0�]` \b:t��F�u�6w-n�*ṋR\UU!;�:������N�^[+/;\�?���>ٻg���U������U�N �`6�TȷR~���#������j�`8 �ۊ1X
I��CR:��%UZҶ� 9 ත�6E�  �X:�hp�ka�5��m��;t�
�۴Թ@�<��͆uKօg��Ư!2�3�
�T���0 Nt����r:m>ee��!����g�M�����,�p��f���@�4�z��B�bB�O�)!+�@8�Pݶ"�w���m�M��e���E<�fUj몕j��V��)k����غUU�S�<�]�Mm�T�F�^��&6�l�ۖ�����ۢ����H[FӦ��v��%�R��
����A�����N&`�T��3���lp�m��UA2�헣�\�۩������ڭ9VX�:%;�SM2@��[T���S�9�[u���U 7`��r���2�u�KЇ5*�U]B�P�V/m�IӒI�ƷZ�kX 
ID��f�A���	-�a� ;N��@[UR��ue [ݶ8 �"@6�Jl	P+m[Gl��U���J�l���V�6˭��L�Q	w3�Em��ydԘ�eyv����u@�Vݴ�b5]Ҁ��pJ��*�>V(`)X�OU6eU@x
�w��)�"튠��a&�ٮ�H�tN�Y�P*���V��UT�H&�
�5kjm�$cEs�Y��6��n� m�m�Zp���+N�����d���R�
��][WK�J��W,pl��;�ib�j���.YI�P媭����7c��������]��2�3Ƃx8������%�9U��cT�ڣ&�<�v�\�RY]U�C'���CІ�@]kl��C�>���Π[cP�g���XgV�Pz۱>S\��ۤ�6Я��t�K�uJ��6��� V�M�V"�Va�f�6��%N�
	��3u��2G���� �wD!t�/UZ]�E��;W<�n�6�*�$��$��y痭�bČ2F0J-һq�6��ܲ�D�y�����-;ci��Rޑ62��E����L�o7�x
��n�HX�-KR�T����YT��`H�h6�  �nn�\ @-�P+~4�UM�0��2���'@Xh0,Ӷ��T�N;�o��?*� �V�U*��4�T��In� �����YD�Sꪁk�*����p��J��PR��@ጝj��ET����mJYA�ܙ�3���ҸH�dm���m�X6��ZW�v\�6��W`9�Y��ښ�.�K�g�ȝe��8�UR��D[n���h�T�����]���5�9�;�r��6���B�)vz9��U����Uu/惉V�C�����Uz�bj �cYf�H �S��^�Ra���-�T�.�sUO$���Z5'C��Ps!2�ck��)P]�Qij���Q�7Xr�*��;uE;6ܶ��rޤ�u��5U*�̛�Ѥz�Rd`*$���j2]M*�)Ee+n�L�����U
�筲��өv��յJ#�K1Β�"�꣗�	��[:�w,����dMʑ����X��=�=�N ڀ��
���@�R��Z�c����|>T����� ���s$�n)[j�B1Y��@Jm���¬+\��V���1������k`#;ﳫ~
����l�۠(���^�"�@烉��L����������p�N���z��__��}??c�W�p> z���@� �j�(�1<�u�Ȃi�`p�hN�4 ��"��J�n��"��?��W�(�B�H��/A
NBX��:��(A�*@#`Q���`&� P���t�Ѧ�<O�DS�ا@� �Q�t I��#HH�C�� |�YE-����h�`#�.�AT 裵�
Z'
|�
 ��]��T���t�u:x�D4!i� ��Avh" R&� ҖZ�Q�W�U�{�D����(8�D6�x��T����
���,���ʆ��кx��ux:]�-��gF�4%���Y-�H[�;s  ���   $ $6Ͱ� hd m�$�@$��i"���  ړ���I	�n��/;6�����D��$E�;N���V�[\,a�T�  �E�Cŋ&�%�&Con
Ȯ�As��C�
��s��6Z��/f9��y�8�뗂�ʪ4e��Rd֚�[;!5�l��9[����ͺ�ֳ@%��Ca&&�#r� eu¶ݳ�k��i�F;yI���m���n������44`�:y�ڸFYZq.���v�4B��c����s�	p/F�SO�"�m�9ǔ�ת�gC-86J�f�v6v�عH�MϢ3�0�s*�jT�J*k:.+�r�Vfn����;S��v�+X��Yr�8q�3n�\��Pܡ�k��/i��O�H�"\���!�]45�ٸ�\�s{eɅ�/���t��"~���ڝh�j�K��<(�''�w��.�Ue){r��:����6�\cc���e{@g�I�٠��Dn^B��+��ѳ�[k��[���z֣GF�K��l=�ټ�[L�/�s�%��ˋ�&5����tPL'I�a�o��h�L^j�?|��]�1�Wi�b�9�{��[���]��n�3�RʧЮ��!ޠ3�E�E��\ =�$G1�Xx�iXЌ�X1
86]����L��wK�2!�#" 7��*��U�"d�<B����Ύ�v��;�~$��Cu�׏��\�u	�B���1��3*���:�	�V(�Vv��:.����g�\|�Os�H��G9X�>�ug1���b.�#i�t�$@{��@� �#����Z�wH�	�T���U�">�vO~�_����v"�F��ڍ�AZ�ñV�
�9�w��3�eC�K�D����!w��Uv݁��z��R!"gV���pn�ޡ"> sE
�RE��ܧ7;d�������f�*8�Uv�Pm�J�(5�<��iyyQ��������#����Z�wH�9�s�@K�J�Ӯ	琑�����]��G1���b7�P��R��� �1��� DN�!������SV�vU+=C��U��5Z�T�Tm;�(|r�ݺ{f㑙��VoO��w>�"��t� ��ƒͮ��q�Jv�j���X��.�����|���֭�D�p˳��f�fO~�����hf 7:����K�E�h{�n�$Fr��՜�;�b�������"�BDs�`}�T����:�b�	8�ܮg�.7\j6�x��:ҥt.�ꝋ�\#�!"1gGB�i��b��X���C���/�T�$@{�H�bx�Wm��w��!����y[t�$G@$�y�����%�)Uw>�Mu�D�u����=�U��;�b�������"H�y�dB�ڵJ��s�@H4D�H���mV�]:��G�BDbΎ�v��;�b�̮O!t��V(ݴ)ۋ��㚲θG�v>wߧw�����!w��Uwwh�!ޣ��b3:��+n�����G1g	�Z�9���"��"!+ H���=�Dm8-.���H�b^�,hU���\`mŧ��}O@2�h��Z9�s��#���T��WN�$Z��Gu��Ю���G�G1�oش��K�Hմs�n�"�S��]��C�G=���w��W�[6u��L�+XWl:���SCP�ŻlF
��^k����m��A�m��]��y�����o!��x���q*���r���טu�2��u�aų���䓮g���v^����n�Wt�N�V.���[tGb=���}�L'�j��!���3w��nK�T�� V�2!rڵJ�]�Q�C+(��T��u�":�1��dB�&�/�3������V�p5P�
���9]��C1�Z[��*U��*E�� ���`,Jl0������1�����;�s��9̉y;�K�D}�%J9�{U��-V=���{G{OL��y/�y�e��rZ�]s���G*7A���?(H�b�j�+ts�Q�C++ho;\I�LB�3�tڸ��-;iͦ�Dhm��KB�
�Zhs_��C�B&b^��3rBJѠ����n��j�CI��!D�?���L�,CxM�A����J��a����	Z5.K��CD�<MC@��\��R/�'�C��p� 8��]���s�6+�l6b���C1y��
][G�S����ُ��zK�]�4K��D�6�A�ӽV�8�]��2!ޣ"YG9������u	R�b��YU��Z�=�r�FD3������*Q�P��F�� j
@�~��B��ʵJ�]�:�b@'U�P��ێ���w�����:v�����u�"<���H��d��Wt�lȇ+�s�F��K~�%J>�#���]V��3�Q�C1�dAy�t�y�<�yA�ш�F	�D������#=��Z�R^����Ʀ�RV����ˉ]]ȸ*k`�ޭ������� �&̑,[Y5��������Ջ�<ώat�f8��1�5ߪ���x[��&ޏmw�v#4 a���&���aԐUaصVw�s�j����i�ipH��P��/1�+t�Z1u�3�Y+��Dy�$@f!���Wt�l�!��`H���χ���.�]���I� )Qͺ���|�d��g�i�h�Q�7YUx�X�E��
  h�H E?Z2!:��43�PYv�>�}�7P�{��]��b�1�]�����"�BDs�U��Ĕ.{u�UڷcK��˒��Um+��C�G1��VEJ�:��i$��!����
���9�I!�b�߱io�.k<��9�!�uZn��C�G1b6��󫰝�É[�W��X�f�lr�O�D}�$@f!�Eq�Sug1���b.�Fӂ����"9�_��+i]�1u���d�p	~��J�:��u	�?.SyWi�Waа�ń,a��xK�XjT*�M�߻=z�f!���([��"�y�d^ +����wFD;�dC+(���yݧO�D}�$GA"U��V�̈w��=��zI'�����
�+sUU
�]���S>��RV�,������of���ȫX
a�K٬��Up�ֶs���;RA,�0_ָ����E80l���y�
,1�,�Ƨ��+v�5[�nV-�b�m�b���@{�MG1�>�m+�`f!ήP�C-/�2
�N�$G�_ I�����R���"���C1�--�R��(��H�b���T��wh�l\�nMl�
�nA�膺>�;�s��9̉W���"D�H5@U@,bCkhȄĨu�U�g1�h@@ T�H���m����琑���+i]�G1��2����9�{M��t\GcQ���Ǉ6�_�\�Wv�\���}�>����H�w�I�I�̋�
�z��H�ȿ�)pJ�y����� �!�i���!ޣ��VQ�dK������1��dFrU�R���-�֞Wvہ�y�sAs{��k�s�F�6�nK�T��!"1�}J�WmQ�C���d�T���'9$�3=�U.���w��̙\�]S��b�V�g���Bh)�#�~����1fB�t��9����d^j��Rw�L��*�a�s���L�si��Z[�����<���Y+�I4��A Eh;	K�(�`��T4�u�i��EaIgd:Y�F���e�1e�7���b�$%m�\+WI��4l�ш���\
F��,h�``�`@��X��Z\]�	f�1��ɛ*�Y5��GF d������Uva�D��������Cv4��e4R"�X�@���������֫Z,e�@�)\�H�Z�5rky� 6�m ��� @��p	  �	   XI��Im�E�'C�  	5�̛4�j�ᡵ��-���]CT���d�R��q�U�n��N�l(]e6�f�<E������Z�3Y���B.���@�@X�1e ��J郒��$��И۷]j(q҆�p�w@�nE1�4 ;l�Z�y���Ԧ�݆&����.ƛj�7�v{\�%-��.����x�
r��-+����-v��۲�������K�� ���6�E�'&qa���.1�c��T�d�ڇ���f� �.m�6��t��f*yw��1Zt���@y�մP�+km�ؓ�I[�3�#�"��GhF�v���$t��q:�Z� ��y�ċ��S�5���M;c<;��][�.Nb��W+mbʖ�hL�6
������N�UX��@��ʀ:R�G�S�l����3UwWuye��w/iDm2�wN�������[��*�\<26�\ȕ��=]]rIl�^J1��x[=qn��&�:�FVi��lwi��͊wYʰƥ3����:K�c�=��=�6	=<u�g�A�Z5���}��I'��n�Wh^�9$��.�sM��������--�q=��n�,��Wn��g;���ߞ����n��f���0�nn��m]��'y$���
�m&g��3?����m�inﻻ���Ԯ������fd�VAj�]I�I3b�кJ����������j�v�V�g{����P��JI�ɘ�*��,��[�!!���;;�k]�u�yNN�I�����L<�w���t*T}�m4x0#�c��Un6�ť$�d�]̮����fw���/��Z��Rs�$��,R�
V���zN�F��@T�(F¢�2�J � (
�E�� �����.��=�=��^��6%��sSfMf$��X��ӱj���g;����E��ӓ��fz���a�s���A�ۂ�H���"�euZJ���332	�(�G|/_�<�eH�-v%t�D��977m����j�퀨avk[N�aIn!�Ꮮa�2�4ms�k{��e�n5��9����u3d,�v���6�(g@��=hB�u�g�<��G@����J�?s��~�Hgx)v��;��f?b��E)'�6�P� ���J�P���c<�^j��0$C�FH�P9B�뫰�{v�ƃ�K�gT&��$���G��C�
 .m&��S;�쒈@�D3�����EMU�\@w�պ�����z-]��7P����>����	[|��'��m|�q� �v��������F�[�I#�$C1���un�2��!�Cu�g���Wn�"� 0	�#@s�_U0�> �ݳ$ch�$V��ԚۥL����$E�8��h�Wj�1"W��o�ݸ�qUn�D�;�$G3�v����/�#��#��1�<(NpR����bP�fp|;!�7X�u �e,`� 'U�x��9Ry��mΡ���Ϫ�Ϳ:�	�V(�V�΃����f������d��Ǩ����	U�]&���c(�ͤ�����?@��BD_�z��j��|5�!"5$c�	�v����#@XEĕ����I'j����Yz��+�5��B5#�ie����:��ڎ�=^�-M��O�彳���Y�ܽ�A���H61��"G3G���P6���W�&Қ1-vnȷL,�e!b&�3%Vr_ĭ���*�>���}�����t�4��� ��R���7WMM��w�(�	�c7�/;v��A'���?}�	�ލ�����y�1�߻�I����. l�XMq�]+��ҽ$һi�t���=@n��No��ee^K��i<Ҽ�6��4�!z��< ��И�Wh�/�|I��3(�X����> �s1�CH"�P��U:vFn�� 
�;�H�`�_Ab\�������B�v��b�Z���r�z�b�P��Վݻ�Guh"��wu�FpJ��Zj�3�|�x�6$�=-B|S^&]%1e�(�`ۺ	�u��Cf���*̩���U�)A
��ޥT��݁(e��~�&�2Li`mc��(`[ADH����%���Q��T@�_ B1(iJюf	~kZ��uK4w���IbƑ��4]E�v�	���L�\��!ʩ�'��:H��U� Q���a�h)+�������[�Q��瀅��z�[`��0
q�(����P��{�o|�~U�J��k>�"���=�L[�y�3�{�߯�Y6�t�z�QhY�X�.��\�
��;�_���e;�^v��">���9�꓿U:vGwY��3�����V�EJ>�!�@�!�< "wv�}�]f^]GȆ����2���ot{έ�uvE݊�ЛM^�*�O�X��n�����ׯ�v�b/�4�j�3�=2��#~��5a�_Q�P�\���o�Bc�к2!|FH�ԣ�Eyڴ�$G��9G1�C�N�	>�ϯ_+�\��s����^�r�]E=p���eM���P�kg
s!m�=�)i쌵�� ��^C-�;2��4�<w�흦�a.-,�b�`���!����'1�MJh�z�$�wI<�b]��J�.c��h&��j�[�݋�H�5�Q�!���^�m���my	�?ĐDC��]�j��!}G�g(匪�n�u��H�s�dE�Zq�t��1���3P�������y��tG��7>���ubݦ-��������И��d}��τ#�,Rs)��[�� > !�c���=�46��IϪ�;!� ����G��E��UyZ�|9GF�챺��z>^����.�]*��AٷS0�`kQ%2o}�u�I�̣�0{�I��"<���9�B�ZzںL��}C�ku�����ݦ-����}���1�WWFD7�gwY�O�o����J8��^ӳ�]M����v�>�}�3�s���݄��3�2!�����һ��<���c7�y��mQ��2F(t�"� (�s�ۦ���G{�fQ�����PUt�@�ͮb��pm2�d�t��3�2i����<���nӺ|;G{������ }~a}?~%��&G��3T������::�[|�#;Gu��vFHƑ�T���n�D��C�T͵��Ҷ�	�x�m�V���8ۮJ��^�8&�l�'%�|G�3���ͱw�@i�s�xC6�]"����F|z�z��9-v΁���'ԏ����	vt�D�;�e��ٸV�	+�y�$Z~J��w�]�j��!}FH�V���Bt�V]6�<���9���.���ī:�W�,	�y��Ǟh��>����@݆�p�: 
(����|���O��A�f#Kv��<Fţ��ۋΆ�;��/|����B.�c��N�̬����E۠T³�f!��vFHϨh?D
�_|��.A�ԭ�|;G�C1ڪ -�g��]�j��!}FH�Q�t+��]�mҤ 8�n�֚5�����$M�}��6��=��9��}M���fH���4 BQ��7Q{��	�j�Q��IQ�Y@F�T��%$I`#�zF/�i���G�p�����5�d���Ev�Z|��? (� P�s�����7��3��:!��i.%�����d�=���ϟ7}�����N%X�G�R���h�f#��h�T�w��v��B���|�Q�9���n�?��d�}��=��D0,��u��W��d�rF? >�E
{G��>��+E?�V��n�7�bxJ�:a�\9G�C1�c��xUں2-(
�������y�]�V�b<���4#1�h�t:7�J*�Psӛw�sGG�����rR��wô~ �}�$FH� ��b_�,4YP��Ry�!W��f�	f�	f�Zc*�`a��.�6�IKM'�QF��`�ib�F=4Rbl��mÀP��ڑ(����Ui�-4y��PfU�F#8���wG`�7(��X�B��c���2��BXA&!-h��¡�Ubܤlr̒f��L ��	�=�aԛ�(3R���n�N	?W�O^��Eh�FT�Yt,�o[�JU�ܜгJ� �m    Cm�H �H m�۰h����h�������  CM�v�^(Eы4��umI�k�u$�uq�U�V�9)�n�Ȑ�it
��+rЃ���	��˫��8Dyճ�W/-��Nw�1�ԅPe7[�MsC�\R�(	�������2[��r��]Շl�@�5�K��AR3&�  p��@j�d;jP7���u��K�٭�i���b��8+�B̚m�;n�}�)��rZk�l���/b�8is�$kv^̇�-�F���ى��v�{q�:|8-�]�d��8�ds�gp�::0���7(=��]�4m��h�B$�&4"��������#�Z�2�躛�3�5h��X��<jE�ݷ5�*��l p��ݮ��Ӱ$��v����[J�T�Z6��e��-
�=8�ʖ	I�b�۵�`mv������ʵYu��*��ۖ�y�jb(p����:�`c��F�-zʵM�VZ�ج!
��������Z',q�A����9�����T��M��5Z��%���egW�n��up<T%l�a]+V�۶�ȅ����hp����˦�pn��y���������?ͫ���ߙ�ߐ�F���6�5W��
[G؆�;���1�Wj�ȇ:����~�)���˫f#D
�r��X��?%����ڶ�7Q�|���C3��݄2G�:A0��i�X�<@����7��nh�z��wÔ{�4R�GwY��y��mQ��/���9yC��M���#��C$��;��Я�̠��Ъ�Ӷ�un�i][J�&��j�fHϨɤ|E��L���;�ôy�3��,}&ed|������� b�`�@� }_����}GF���ڶ�?o��c2����������	���Q��{�]�U!t��6*�6�âK�\�fm�Į��{�ޡ���Q4��߾Q+�mQ��/��<�����!�}ϡ痕wsG�S�rߣ���r������>c��}o���$��g��R�N���u�s1�ϽSlgHשE�f�`��ү���bB+{4h�/+#��ot����=;���V]��k�|���BA�wY���!�p~.d����f#~��Yw����D�"�
�=��O���>^j��tdC�FH�Dz!�������W�k	��m�5USf��r�7ji-����0-R����qx�riJ�L�	�1��cغ�l�%KNYe�z���MJm\It���� �6�tε�F�쪮+�� z(?*��0(AV)R���t��z�ø�ɠvXDttq�n�L]�n�n�>�y�3��� 
��L��.�1ns��S�� ,��(H��!�����_;T���� �FH�xQ�\���~�X(���}O�}o�#���ڶ�$G�?h	'�#��f�_�W�� J��f6W6��7v�a�wIR2F}�dBDoOPYy���+H�Q@�O�@b8{�n���y���Z�m�"� ��4-��~��{���n�>�w�Ȍ���R�v�2F>'�@� Q)��>�ß�z��v���۰�(wV����WJ�+�j����!��CwX��O��9���9 $�����<�Ϳ�S���g/+*�y�;�/j������G���*?k����#��F�<�7V��u�?D��>�����G��m7��ȃlհs]D]$���[V��hȇz����=��Ww48�N�<� %��6��<�M㛯�۴��3�!�$��Cu�U�MU�>�N�G�Qb�1V�6!� �RF'DeS�V�D4�� M�g���w����z�>���ٗ��kٌʺ�wwB�bݫO�D{�3"2!8�լbUJx���NX! �8�<�G��C�~�����wQ���FH�2/5k2�����@�������ﾷ��{|������y C��*@�9��y�������8���T\C��Ut����\8"�/.�v^�����S�[{6ޘ.�k���<��dù{e6)�9��k.9ݙ�(�rntsW{e�NLfN�^��v�>���`Lmv�S$j�wn�Wi3;	�A�R�O�q\�� �X"Y�h��<�͜�?=T�գ"��"�u��to��]���D�� ����yo�S��w�j�H�� �b;�n�9�S��A7l85�fca2�&�f]���$�HH�����˼�?}O9G�W����jƭ]���H� 6:����� �R�{�v�u4}�:�-��|�&j���d�?�S�@BE)����f����#�N�N��>����}�Gj3e�S��S�;]�,eU�Ur�?(���F��ys)���n��ߙ� ���W�">��I+�u��ES��[�Q��	�U0� �-�@h ���� e�#v�#��D< T�r�!�!��PQH�D�S.�Q��^`�)�EPT@��Ѣ�=;,1�]�F96F0�5B0Mcw�P�$
! D���.�)�i��TU-4�YQ����NG��j�W��偟��/���P8�D"hSG� �>D0<�D�u�܂y�����G�BD?��A4
����(����?|���gwY�G 0z�{S�5�<[�mvI���2ed0�˩��i��o����}G�|��:��g�g�FD$F�;IK����Ē>_|��|��=T�գ��s����!�h��p��Æ\�yO�?{��?/~~Y�|ߙ�����%�%B��wL�a�e]�������'��i���H����;���ך�v�FD9�? ���hhWmW A��>�ϲ3������
j#=�3��~�������ÖTg�t�bWAZ�t���+n���!h�R�����F��^��׎��m��f�B�7�ܙ���Y����8�%2Є4[M�E�س��t�$<����㈙����u�l4��'�w�I�S��ϑ�ߑ�1: c��d_��#���߁�?�[����}�3��ȆT�黲��3�#";��`ܦ-�|;���H���`}m����T�V^�in��Fꝋ
Һ�wWm4dC�FI������?�J��j�?~W���2#،�9T�ZVd���~#�� ��������$�
v�����H���聏
v�#"��� ��w�?�~���~ַ*�Lʶ�apʙ&XT%阚ZƆ	c3>O���^����g4q3���a�s��EP呂H��!����>�1m;�yx~�D�A��QL � �QE!T�E�iUs�iמ���^L�����D�$-�������Fw���j�$G��2#"�5;U׬���Ъ�M�Vw[��`gj�I�w�;�����V~�ϼ���H���$�t�dG�BDg�_��}J����$���~��n��|̈�:���Ā�g3�CO\�-P��e�F0i4Б��E#��`!�F�e�
����8 ���G�^�s1�}��=�+�+�?,�������>�[�cVl��Ҷ�,P��m�t���ڻ�y	����mc���Gu|@~�	؏�|��/���>	�bDo�fDdFs�U;V��$>4}��ȏ�!����ԔwO�D{�$G$c�I�:�MRN»���m�|���t11��]���i*fތuk�3�K�ش�f��b͋f�`�YSf"�MMű ���0 �*:]�����W�]-��e��і���p���g@r۶��ժW��J�|�H�Σ��ȍ�C�W�"=���ʝ�P�t<qŻmG(ET��<��4�';]L]����y	�38g��m�dCA �I9�~��~��}��\�e���G3
s���h3j��b�t,+���D}�3���;v��#�G@$   �~4*�>�<�O���u%�
�dG�W!3�s�ٝL���LQ�H ?ߐȏ�ߙ����_���fDd]~�𿃬]�<��3��8��������n�$d�����	��O�h (����}���a[�|?�#�!"2Fo(O]��hȇ:��l��P�HF�L�)X]�%�j�0(��,�ϕ��y��-ߔ����̺�=�O9�2#"2�,S�iY�1��H�� �5ߐ��  ��ޥ�����;.�$Պ�fM�u�
�X�����޾��FH���Pv�ёi���gua?B Y�''���hs�:뵼�OQ��V�FH�|��a'�$�@��ß`�L[���G�BDd�eqE�胢%����	Ynְ�(л��ёu#2#/���j�$Z �(I��~���X�jҳ$g�C���Cuڝih�
�> �_|���wu����U�"�2Fd@�,D�E6�"�e�r�(!V�	��:
Q����uI�X:�ѡJ�4��BF�6p9���Sc�1l��9dqJℤ�捬� �5-c�[nHt0�d��y+������A��x��5;ǧ]:�i,90 @�   6�`  ��m�� �[R�Ӓ�)�  @��ی�fX]SEҚ�ҩ�Ur���\�ne�Z�謔��5�Xz�84<s[N��r�X���bV3�Tr�i邭V�WRI�z#�U6U��v��9��-�Z�j��T�����(��D���1]&筛r���Q����y��nKPX�z���C���;o<XB�I�a��t8����b۴�p��O��-��7	��bź�>�l]���KU1���g1D�6ym�Vr�zwvsZ�����������[rv\ڹ�83[k���4�@��p�졉��'n3�oR�ު�,L���Ł�mܴ!��m����Raxe�3uJ�l\:�C�O�-��sݡ������%c-�jjc�\54��̤i?���{�����h� �C`iMgJ�u�w6��(	x��{mw8�I��gZ쩰Vt�H;���MU��g�#�������n�D�V�m��Ldy6Mh�X(��ᝎF�<�X���J�V�����$��]G��F�ˮ���{7b�iv-��w���fE� 
�J��U[�	�g�FD$_���Ż���G�_��GwY�C}vi���:�����Ё]�\#�y���ȩ�.�)з4�1�a6���>s�)ڴ���=�;�@n�ͩ���f�}���2	@��Sv��y���]<zZ;�s������_���bT�"S�V�FHƀ�Q�Cu��/
	�e��i��6���6cV�W�}�w�?�$FH��	��7FE�]�;�����7�zVe�����Xq B[��;����)ڴ�z�u�VQ�C �@}g�V�K�|W��w�H��c�v(\��KNvnF1��q�,�񬏞W�H&�v$�H���dA=�e� �&�=�}��/I�$�{�����$��<��$�}_KA$O���$�{_o���n�$�H���A$��bH���}�%�$�ĐI^�S��*]�7�W��X�	"w���O}�D)F��`�D�ܴ�$�N{�2���h$�H��%�$]�ĐI9ͦA$��X�	"xr~������Q�i���jԌ��i7�O}�A$M����Ok�i�B��'�R\A'���}���В	"}�֙�N�e� �'��\A=��I�5���U�eeV�pI��X�	"m�%�d9�A$L�6��H&��.e��	 �&sIpI�k�$D�si�$�Ȥ���$D���/˙����H'�]� �&��i�$�f�,I�3�K�H'� �h��H��d���@�!��!m�"T�%%��߽�(�2����WU��|����.r&؃������9;W���kh�w&Bq���Ic4���8Gp���kqӆ�[nx�bM���;+��y:Yk�T5l�'wu�7�����D�IFT���!��}��s㭒��˭	 �'��ZdA9]�$�H����	�݉ �&��L�0T��5�H&k2ĐI}�.	 ��ؒ	"g9��N�H���8�.]�ք�I�.	 ��ؒ+��Q?~�i�I�}V$�H�s���f]M&��	��bH$���� �	=��I�=����	=߶K�e]愐I9ͦ ����A$L���N�>m:�>�z��7�-
e��WS�mc�����:z'@g5bH$�����L��I�=��L�H&�_�L�	 �'��\8 ��1Bڰ����"!�T�]� �'��� �	>��S��H��}�~�+I�$�}�ؒ	"w���$�O��A$O=��$�y^���BH$���dA&�Չ �&sIpI�nĐI򧽘T��n	 ��jĐI�H��L�H'�]� �'�}i�I��n���TQ�6Kk2���Y�]����'@�����"k�ؒ	"g9��A&sV$�H�s|��fYZM�$�nĐI|� �	3��$D�i.+�*�t��K�e]愐Iﾴ�$�N��I��P"TT�HV&РT�K"}�%�$^݉ �&r{\�~d�ZM�$��=�,I�<���	��bH$���ZdA6xp��r�$�H��IpI�A�rĐIﾴ�$�}�ؒ	"~��eoзt�)��������hc(�/�6��H'�]� �';�L�H'�]�ʰj	"}�%�$���%e�ZA$O���!�0 �|�����;�3�j}مJ�&��	�݉ �&��\A3��$D�si�$�i\T���w.�A$L���	��bH$����I�]��j?�,��X�	"o�;�fYZM�$��$D�;i�I��V$�H��IpI��Z������c�ۗ�Gl�i�BH]3ګ.�6$�H�}��A$w�bH$��ԗ�O}�A$L���R�ɒ���H$�ڱ?1�$�甗�O��A$O��� �	���/+*�$�H��%�$]�ĐI9ͦ �	=��I�7�=��/	4��H'�݉ �'{�L�H$�ڱ$C�D��K�H'��zJ��.�$�H�}�� �	7ެI�3�K�H&sv I))ў�˽����r��]�N��ldb�j���S�GW[j��ە�=l���{]q�4�wc�v���Ӏ:�C��'�7���M�����59�eH�����1��X�����u�&qYb�su�.���t??.�$���\A<��I�=��L�H&��3���A$L���P�';v$�H�}��A$}�X��	T$�ϧ;�eI�$�}�ؒ	"w���$�O��A$O}��$�Ou���WY�$D��m2	 ���A$O}��$���}�X�	"kϧj_�+*���H$��$D�i.	 ��ؒ	"g9��A5��ҳtL�'up9�k��&-s�ayS+BH$�ﴗ�M��I�3��b	 �9�A$Mu�5sr�I��A=��}�Ź�=�m2	 �U� �'�R\Oʃ��W�t���]hI�>��L�H$�jĐI=).	 ��ؒ	"c<��b��I�$�O}�A$Nv���	�bH��ﾴ�$�n���/.���BH$��ԗ�M��I�=��L�H$�ڱ$D�=;ۙl��H��ˠj���Uk�B�<�� ��ؒ	"o����H$�jĐI9��$�L�%틫�h$�H���L�����*ĐI�.	 �}v$�H���ʗ�J˽&��	=��I�9�K�sP����8�	�ᑎ)T��&��Ӛa��n��Pz^���!x`���q�F΃ZM4J	P��Fw(7�w�]A�LY�j�'�`T%�ȅ��D�Z;4�3a���7I��.�E/C�#�<1�$<n�|�G��zBS(%�����4�$RrI�"�`��4kFo�����6�mC�D�z�0�������v�Qm@_ڠX��חbH$��{i�I�L�ʙZA$N3IpI�k�$D�si�$��E���A$No���4��H'�]� �'y�L�H$�ڱ$D��K�H'� 7��j�FJ���`X�9��4&�uR�]��kbH$���ZdA';V$�H�}IpI�۱$D׾���e��pI��X�*	"q�%�$�K�$D��2	 ��h���Wwu�$D�i.	 ��v$�H��m1�I�Չ �&v5�fUbI�k�L��I�;��dA'�Չ"@c���ԗ�I�s�&ee�hI�>��L�H���y�X�	"}�%�$�����t������T�ٮ�M3,vr�3��R:J��OD�L�I�6ޒ��	�݉ �&s�LA$;1��LV�H$���\:r��7��I�9�LA$s�X�	"k�<����4M`�	�݉ �&��i�$�L�I�3�K�H'���J��.�$�H���A$s�bH$�ﴗ�>�}�$�J#�h�SӾ�U+�"�b���	�
	E4��禬�u�%��U[,tr�7jk0�
�"��&`+g.޻�����]��k<(���.u���;h�wf{M,<p*Y�r`�s�.����Y���H�-���_<5�.:0K�U�A��ӌ�� �GS"�{�Q̌Ȍ��jRWU\#����o�
(}�}b�յg�g�G���Ҵ�dG�BDd�rT�V��~!��i�����S��S��2J���j�^X7V`�������}�{���!��Cu	[�
V톎� �	��v���?����>�U�����@"�~GwX��o���`n�Σ$bD%s�)+��	�� T�����Cn�s�M!k��.�n�+�˰�ۺ��mY�1� $BDoÒ�ˤ�����7Q���Խ��*�����h�а���$l}	�]��Z��u�����f1��
�Ck}�JݷH���D$G@���tؠ��Z����
If˪�I��z��j:�����!���A����7��07P�Q�1"ts�)+��	�|���}�������];?}��D013�v��.�O�D|����*�Gi�V�a9o��F�6�[i�8���h����Q��H�x;5�">"w�����#�D$F��U�w������Cu�c��vӤ��	�2�bD@���hRWv�i�wwuvz����Ѩj�B�ڮ'r�/����I��[��VCvF�`�n4>��<��oI(\v���L�H�f8�)X�$�g�SGRwE	v�^��8�4�b��[I;åut��WD���bD4�(n�8��]��gf�� $BDoܨ�ˤ����!"2F,d�Uwt���#@�`w���f�7Q��Ĉ	r�m��-�bMc,B�Z��J��'n��d�{�	��'������_1�B 'E <�G��o����Ho�[����# 9+���ꫂD}�1":n�8��]��gwX�!"7�P��	U۪�A�a)�p�0��9��ɚ�?;�ӻ�BE�!c ~�����s��F$C�>7�~������� ��_U�d�j��L4s#�D>#u�`��B�w�������;���漩�N�	kl�+A���X�Uk���u# 9+��I]UpH���$@H��]O��������B��>��+���WW��7�<�P1� 
 
Kb�@�UWwL	�Q�1>�����q�af ��t0r�*J�M�������bD4��Bo�);�a���{�	���U��D������OZ�I�"�2F>�;��j	]Upn�=�1"D2�˄t!#�b��儩/�Ad1�J|������ Ab��I�P�"�"T��"F#E%5ڞ]B�̙@ۦp�df�-��4�5|Լ廀  $    !��-� [C m� 	� :Am-�l��  �7o<�u��ĵ#�m�\nI�on��F.R�W1v����KB� cg�6xb��nVݨ8:ca���{Ɉ�)��7aonL�k����R���l�a� �*�6y���v�`�K�r۷ma���ۭ��8��U�M����udO&�6}Y�*�6�.�ى��(i�h��]���&yi0�up;Fe��P܁�R$-u�-�@^S�Us=�[ڞ�mu���2]W��1E�&���N̜�Q�ɰ�e�V��5��ӢZ]�������N���n�x�{i��c��)�sy���ր7 ueu<��r��1����W�2B]�,]#�B�������(),R��H��9.�wig�7`�!��aW.���ٺ����wԓ�;��@�O@�x��1`��3�wwi'���{��&�n�:eQZª�Vz�*hj^ŻlF
��9��� l�*��X
�מ��G��rIk��n���&���us���R�m8�jާ��<!6��<�Y�*z�xk[�aEL˒�/$,��3�2�ֲ0�{�����?�j#w�P9t�| ;�$FH�@�UWwL	�Q�1"�cU������bD�d�j��L4d�~�s�|�{���ϩb[����B�d��j�7n��;���w�"�BE��c�����`n�Σ2>Ԉh����J꫃u{�n�$FT����vd�{�	���I��"�BDd�J�Q�;~GO^���9�8���Rv����s��� �cU�VW���bD�@���Rv醎��#�
�B$c!2A�T �@B4i�,�A��F�$�Um]�H����#�,S�L	� �gw\�����>��i�,�&"�˸��J��j�]'h%uU�">���"0T���V����!"7x"�.�o�D|���������s��ā�%hh��0	�.4THB�4,+��[G@�sݖ�;+�D}�1"DF���Q�p���N$���ꓷL4d�{�	?���<�}��][��@w�H���r
�)�&�s�|@��n�9����WU\���bD��R��I[�$c�@H������AED�I	8�I{{�����՛*�Iz�:�K���s"�ieĮ�[��LKR��Иz�U�A��<��sr�w8Ĉ��uv�ӟ
��Z��e.�z�k���k���z������m�<�n���m��A���[~���H���tM����@ W|��{��N���w�H�����醌��y"#x'e%WV�$@i#���;���>_�� 褼"�m��8��XI;�b��wI�"�2F$@rW{��My]Ex�Q;�Y��<�WWi+vd�{���7Q��B{t���|��̌s ~��t��u#.���}����T�F���b�Z�����J��'epH���$@H����醎HǼ��	�hsw�[Um>�|�`0( �En�$c���b��`H�:���+�������$�X�@n���`�
�ʫwv�*���WG0W��ae����>i��d�������ҥ| =�$FH�2ꪱwL	�P�Hؑ��e�N®	�yg�S˝ʦT(<�5��Kn�HǼ��	��<��.�Iμ;�V�
�zSB���#$c����wI�"�2F$@<�v%J�W���bD��R��I[�$c�@H�����9t�pH��P�Óߧ�~�{CUlQ�G/#�QM�Q��SN�Y��7<�Wm�/6ޜ�H�Q+�M]te���\5�<j&���	X#��4�Sj����&V�ck�����g���<��u�Ksnֳ ���'��M6���Q6#f@b�O��<�{���x��oe���\#�"1|A$Ԟ�S�Z2!ޠ$C1�艥i�H��P��.��J�03�Q�C1̕U��ӫ�K{x��狙�P��:�V�]�8��yr���Uj�b���R�"�-#|��F�M�O
�2�\ ;�$G1�ڴ��3��*D;�dBD��Xi�U�"<� 3~\6�-؂ȢQZ��]��	�4}�w��3~�4�>	�#�����)]&b�@�C���Q�� �ZQR� !kEmR�� ���hFf�$��ĎˌFB�ZRC ��Ae(ă�� Y �$�4-�����,N
TD��Ƭ����ňĔ��B�B,X0 �-��Y�kCl���%Ȍ��t�L�C��F�8�fja��"<���Ί}@=0_F�6(���h�@�
C�$�����sG����h��H��G9K)��Z���z��C1�P��׃S���ݙ�k�yӹ��uI�ҥ�"�BDs�`}�I]�1u�=���Ӱ��D}�$@gh�u�.�.���n���lA-��)(��+�w�:r��*�w��BDs�
k���N����7wa��30s��,XV�'�vy����1"ewk)+B�7Q�P���@�9JS^ufD9��f"��Br�R��ޡ"9�^`}�IX�b�9�f ���}�o�O2*3�V�����r�������5Xg�ȁ�u3ِz���+tTg�^��f!wc8Ca���q�u�q�E�zAdW��8ҭ͓#����d�e ��t0�7e-.�]�i�U�">� 3��j�Vh�!ޠ3�Z �yѻM+O�u��Q��+���u�3��^��
��u	��s�t�UvP�mS�����{sZ��Ҧ��~��ꁙ�H��6���t�7P�	�Gh ���I�@��<��>r���ZJ��s��!���oe���\#�"1gGBj��;�b��\�]`t]��ڀ��k\�͖t'j�i�H��P��.�0+���C�G1���RV�pH�:���
�@�	I$����!�L5A�Q�R뢮���P�f"�ҩ�t�pH��P��r�cB�l[UU�N��Ӳ�b��X�s��ҩd���=^����vXi�U�"�@43�n�$^ �+'��j��P!����zۦ�<����zj!ȄI	ͨ��@�B�LD;�s�@z�j��n�%	��sS5�[*�X%��JЮ	�P����Hc��g1���b.�#j]].	�#���:�J��EH����H��oe���\#�� H����Wm5h'wm�ľ��M��������+�ձ�1l�3n}��.z5��m�
��vzNb[J!E��[LiT�ɨ`���f�����h����$���yc
�oZk6�4+�5��ң�	r��?G|� f!�����n��u��!��s���;D;�dC1���+B�>�g�Cu"9t�Ю��!Π3�G�]J3󃢧ͷl����5=*E�ڻ���"�BDs���V�X�b� �0	�G��q~��4�*��u	�{8:Vhh�C�@H���2����>	�#����ۤꂭ�6R�L����F[r1
�1��38�z��+�Dy�$@f#�H`}
��b�0�	AB,�BSH�
(P��jU�������]].���!���^`}�T�Z1ub�uX5	V�V��A7�oT���<�o���y�$@f!���Wm0��-���H������u	�B���Uv�� T�{�ȇY �A@�y�H;~ӫ$���Ȏ�;�7P!��B�Ӻ�m��4�q�me^V��,�!]Y�C�@f!�����.���i$P�!����\�?U�V-"�2!���j�M;
�$G�BDt�5":<�՗OQ���8�S������<�!碣P��BR�(,���U����D_�N�ix��j��aG�*�\3�ɡ�DQSD�֔D�
8���B QT� K�(�2
���������Bh�<��1��9��Ȓq�gZ�'�4�c�c��S���5�n�C�?�^U�4_Me>��J5��?�{�R�QL6�C��I��N�9�$�*�����?�G˧�ٺq���j}�܈�a;��?_ƈ����GF���۵�|�����ɮ5��y�-����=�R�+�~i�k���_��(//���`O)�s�}�h�=[�O��
[Ett"��,�2Mɯ]\1��H����~7�	�v�z�]�~�x�=]����OU� ��ⱚAY�v&�� �OUa4*��7��C@+ T $AP��`@�BE�B(@*D@$Q0B,AP�P�T"�B$@T$@T!T! T D	 T!X(�C��l]���-8�U��Ǐ�in�{�X�z�$��(.��=��;:x;��{N�������
?Ϡ:=��v�vw&��|Hu%{:ϬOG�{��y�H��T� E���Qc�������Ө�R���<hz�S��r}5YԿH�4�5���L{>>���ձ��6���Y���Z��{<��;�6[�����ٟ��v���(/�b�D���������=�}�=5I�~Τ���xD!�8��-~���{gY�C�-O�ꇝ,��Q�1?Ǒ�Th� u�F���R"(.�0��d�t��,��L���T��Ƥ?��c�9�((���$a�h5u!T�N�]:g�h.-JB�_�`�M�B%
���q����%y�}����У�<⠠�A�z�<1���͡�WhȘ���?�ݧf������r{N<�x����I�&�i��{��@����~������߷Ͷ�>�*
]./�t<C��|��?�`B�C�����T���4�SK:�}��A<�÷�"�{�;7':��W,]x��zt����j;C�<{��5�D����Cd�vgQp�Θ7�������Ta��g^�u]�}er�U��c�<�N&��\�Rd�3�T�9Mx�a�����W͠=ǟ����AE�~��I`{H	�>O��_����~)��A������a4�x��{}�q7�5�!����xx��*퇸�tY�=�t?�]��BA_(�p